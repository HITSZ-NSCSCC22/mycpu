`include "core_config.sv"
`include "core_types.sv"

module reorder_buffer
    import core_config::*;
    import core_types::*;
(
    input logic clk,
    input logic rst
);

endmodule

module moduleName (
    input wire clk
);

endmodule

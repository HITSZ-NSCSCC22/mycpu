`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZL/h6ISCDZfE/v2gfumQecI1Lu0hBKVNHYWa/5t45/MWFxAX8xOtWf/3N8O/3K2oLLYcUWD1oZpj
Qwi2QHM5TQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XTWPgVsVSvOPR59ARLH99gGkhxe2HFkP+Rudj7uP+Rh2Q0hMoWx9LIN1KM/rn51JYIlSe0sWwqUt
TM3Bi5jpXAlUaoHXpW9ipuc+W4+gt5dNJJhlNDZjmHDmmuXz2ptx+5YubxYzLwuXBL9i4paVtgWG
tiEyXSOv01WP8quUMVg=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z7wLbViUaVPr5QNi1P5jvaf3zQ4Y63BHxaOrSNzPHnjUAJg3Bwq8AvQa6bh5afoJwucfoKDMDVdo
BasmKoAvPJ4Hg5KJ/xM2g3INMV9+luCZMGFsfRUouC7/o8RkjMvYKx2IMPnA1qSX8R5uy8mGMBAB
k66jnn0k8t/q7Radx8dI6gLm4zEi4ytcbRD8ft3nqmkIC6jVnoGqIYFzESGyJgYChpdiD3OpDuCM
4QqZAxSXvJ+g0/MnuXIKU3WNEXpo8Y/vLz9DBDj4rjQN6yLghSdkScNmLqol+ZIs/PCEuWx4LjHQ
iRY0Wmxdg71SXvFvoXsL9Cx2JQoB9n/gO8nGgA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kRJXp7E0H9ROdDeAeu4GvNvyIcqzJC/O3Db6ufOENpIzDFCzCX3VfivQr9pK3PPhgxjzMGbG3rAt
dzN+iIMxglVKEyw0FdpiGV0B/F0zyh/s8zyQoBWVWqn0H5YRAzPRXtXpo2fNCj+WnkEOC4ufCHsY
iCP9OCcdUUwaTqZxFMnc8LsptlkDHBHZTK6AXmrnpvAae8Er8rNb0SDlISaWwlwVAefNefHEbL5u
6ii0HW7uHABmKXQhGEVveWYW8pPgm+jdym7MbtZGio2pG/qCkkNBX/+d9MVTlPfTe1UJC2ow6LrC
NRCEY9jryf8l2Xy5rGBCMbi/MDL0NMc7Q5kkGQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JwvOsgNIVg2tH/Yqqj/XZ885o5PaoG/9gp1i8pkh2wWYcW53TymM+JlxACVqFuUJk1o2EfC8Xdd2
mF92i+rpKyVDOpuF6f0u916rx25rV12LW1J6sIFMST3CgHr1ihl/I3/5w5ZtaEWB1Kaqbs2F+wyY
wl96vJc8hY8qOUNWFm4muMCH6PPXNYf7WiqvidIVy8THVegbu148ZTfs1jNUTVpc0uvYXC6h858q
d7lbqpC1bqpe+kgYarCD1Ps1IShALrBd1gMOaHs05AVsIuIRWxef1qlC9scRLNtx167yoZQ9ynSq
A7bHBsga1/dJvFYsDUcEI6Sx0nZbngWQJM3agQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OQHE9sNaN9EGVTcqFQcNtzfDDcbMNEEAVPhJfihF2sXZhfTAiWZp441grlejPi555jQGIbqPKwAW
sH53S/TU8s1hmv6CL2n5Y+9g2XJqD3eRutqBL+PKRINPIIgC+O0EHMrvVrofTVmYVkq794cChXr7
e9KaMpIg2z4JBRU8hnQ=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fvyid14mFMAi+qpMT/T79jmEJ5rS8XliJ2hBb+iLiwHHbVyfVqndj5FshCUyeIOdaa/XjdT3E6rI
kxQthivhDt8cpB8VGb8EVjr14KLOvdeiun4z+MEGe82sTc0bOz2C4H9h/mKgst8Mjcqwts9mnsjY
TsiAYfytsXrj9MUR3ahb7SzAtrUNECCrfqfu9zOtorgX8EPw8N8ZOYautWalrmb5xW7ejT0hYUzI
MzTgeEGTiWlW/ZG01uWD2zyeOV50dpyUYgymm1Glnm6JN2E/to1+u06ggFZI9Mlhr9d3kS6B48kp
T99r5uQgZaiAhZ+VvXv+4dg6BNeL1WXESIE6XQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64128)
`protect data_block
4L2hVQe0/Pnp2a2yE+4VjdGRX6kb8h9FmaVHBJTuU1c2wK+zGXFYYlh0OBEFxXHneIxb/ma+2+iH
iw2uJ4uG6zV2VFkO8AoSoXf6g19GKNuYvwQTWRjBcyEGCyfBGDMRQVD2T6Myk+82k0peIeAXIoIR
DyAmwfJk/MKdUjsnu66TujWieRU1xC3GLuU+vHvgpIq59xgN4vDfHBojeuzgNhZWE/sKWrI7UFp7
QSDK2ynMIEfOzkzL/zejp0k3VEht8Se8LyhBsgNCXCWF6KOQvEw/iCL6jax6xPOWXNO78WanZaDK
7dHiM8M5HFMSpKwlUc9IIRbc43rNWrwVZxyfkty/UWfoax1qHJJt7VaY7crgM2D2/w1CMSy2nc4p
AI69wlpxgF6/yrJlVzx6pb+BEmR0pGlfF4YSjfN2JUXuxL1INhnTd3Kan3zbycIZNOCFkyzelhlu
6l/GFqW30l+KAlPSqN/Ba3zU3HD81AdxG6D2UavfHmsWZtED4m9hiGS54MfrwEgKzYMWVeYu/pZ1
rD6nGItWPhVDtdSLcx76tZb68qYcnoND/nZJL8vRJFmvDA9pWpWzN1NW/8zA3IiAdvET6kAkKVZ9
hYocYQKnD7uTSRzE5IjiNxRfWJbrrmWVBFkoX21mhkmUvbn2j0tWOUS2UasLk0WezAFp9h01acnf
Ybug84EIxqi67DATMGKnZ4R7Aq5qQh1OPIweVsifFeLqGGJagHR77AshtrJmskKhrd+66ST3w/5e
ntHz+sdkeRCqmqWtCP7iov0HgfC91U7E9iEUJtBwVBahMCAd5pNak17UaKoycMISZwmslgS1aU43
54QvNwG3bTy7OPhU3HCIGgvJRMifPS3PCkcJ067v+1fsOBu/73iOeCkChfYXHqrCkfgc15GFzJ5e
ubdpP9MsJqp5m6usZxmHJTSTWlIvGCEeX6Jx6P72kK95+2m4ntSgzsyVkuGScXoHUjiQmgW5g/WJ
SnfjISXg1Env9SXbiOJ2t6CVB3XozrHENpJyK8b365468YQNwpc31vPY3BhqxM61YyfrZD/Ou3In
T34cAB2hyQDuV7JjAeQk+wU5vuub0I5pVkxUwII+D8GBaocrcIHqFwVeFOLW26f7YeZkmfJd8p3c
JaNth3MoDlkYH9J5tHV7k7yjNkxeqlv1UBflj0WoUiNs0tKpApn4IccDdzc0OPIibocELzpZKhSI
geUvqXz+l6ojUVx2Rf9yUQRfcbkR6fgCeisl1CRRZi1LiVebNfJu7bvxdr5g6NFrY+sVtFLoMlGd
4oCGxBMnpOuipQKvix2zqm6hn2JSsQZyXRWSHiV2w9ghCoO0UtEb0Eu9AHgClI271vILwVqDHRjq
qwOFkzWUfqJmhHRVjbije39cWBrZhzvjsYpCa4arI6YK3iI1WESn6Vkdw4BodML8rzbG0QTFfGmn
tfIsnW7CKb8QXhxZqY2wSySDgXqL2wZ8BQhn7W7evCJkwP0zF2Ht68cts42oAcNKy6XQuCDLs6CZ
dZ61iwOmmvL09W2P1bvqCX5qWFIC9WMcQXHwhnSAg3U27ZkCrxNcqCpMOYJj+gIWA3xUvm8drZRY
7zlpg7ysfWwEr2W1Zepv4aK8EV24FAC2c9egFOhAEf59YFXqTSOd/PbNhVEpoVidT524s2HWgjy4
cTIpAQWk+xmdPejPqebm6tOe91eZB/S9FCghhjSPkceoQbYQaTiJPbtkZwXiUn4y6FxlAE+U9dFs
P1Q2APgCG0zttMTfJU7f2t50LDYakLpIgGxgp7zYhXR6X5BmFJpnMulWFcV6gwQJPyM0d812Xzqm
SEef2IKKUT2ekT2Tzthu9c3xhGRLi9/wgetdKu6AXOvPnRlVZJ7eePFBq6FQEcf1oCtsJV3DXjD3
PEBJcpDohQVl68nHONHA7Fdsx3BuhXwJd5MVUxe6j+d8eIydCpAgrGmIvLKg8Ui/JRck/5RWEzC8
oqEEl8ypA0BfnHX0I0XC8uLzll3Tuy+FGK7pVqiVpZMo85bAwVl3t5LG9zt/s/UUcJaOs4rhzWDS
TiiKUHI0Gaf7yqgFammpQITCmOvGLU26xFOMjDbzc+GZ5w4Bg3kawhpRwmDlL2PbPp/joxJ4+iVO
mX3hcoss4R40foaTCgCuiNdvNytjlBnPEdvF4t0Lx0xrnhcY5awSqKLBKp9sa3okFk51hhh7mfVa
4bNh+lkwRd8G9K/MAK5+G6Xbn6klaYWbKE1g9SSVbQRN+qtjgbytbhAZ/8TBs7rDkDFiBghcs1am
WBJa1A/9X7/a3HqDdsAA68zs7P9OQEfmmLJTxhyjFOUaJZPCIBFYt/OCoUBBccWkbxEPf0cCiSVR
+1977RDly/l72/xyX333uoRxs1qLcrybp/yyCYOO/+GK9F7SLyvzVKHv4ZiazhhEb1KSQma6/bci
pnweDF0xweU1S2IIZK+hVD9fAKZyjLMhfrddKbmP+xUwzgoyPDxWZemTRrlJttXDElK9ukY2hOiV
DYGsv6MViOXwdz177NOtSNHIbi3c4lq94+11nTLCy/MM+lCEiOKlj4OcVKLVdI3pxfTkTSiurjCg
ECoWiadAYLiTexHN2MCvGt4HOvkQRDBKUkESKIGx40Y4IAIunH2gPw2n1aTnREQpyzlLa8M/7yAQ
7TSTKEkvAjwS3G8f//Y+KcYNpUku8CmR0rxL3oSkW3rgRIVMoeZbCA9hN1/H/sqqVANOEoijzLVz
tqSml0Kk61mLsHKzHbaO/oIU5+rZ+p8R2DgH9eHOHeHqSXI4GlLCPs7J1eGH/d2h+rs5tLOSxqIq
XGq4NsGQz+q73GIs+PX0vUvupl7hYnAV5Dc5HxUaEbHMdSX0jyJhdZnDQrR9YFFDqfN9R/BXjVvM
VspX5BROVRu0Z/3AICPFQx666sgsPOBstbszbDRaXcHmEZx8T3HMh4fXSnPyAhwCZsG03CTc6wBH
BrTjPLnao429IJMUFYlPjMO0vW9+j0RkYoatkvsxmm5ScaVUr2u+5Bk9GG7sHedkmNOfH4X3ZqRF
+A5GMJGdvnKWOGA6icBJiEvsr0TytduMHPViq92TLg+0q4zTdurgO3EiCWdRynXjhTkkEaHEmhLh
gYTITTsBBjCjsA95yOVXICNn8DBKOnjbUxxNtzpEgx5Jintou0shmiRFOkESLP1yp/41oeeVzI/K
pAu9f32KXa/Hbrm2OpEu6j8huruI4vlsP3b1eTSHPwddug80oUfZ6lkc6wEiyreIXUFnjBwiHKuy
Wp2Lp4NFpKrInlV/T9DStMrj0Lr3F8H5sT0mg6vo9NXUxaoSJpaZTXIqQkBmpGVNDhzfHnDKLkvB
32ro+dN330UahxaaNDustXGlUczDwLdVmi4dAacRKjdWOssgtyk1i2SsVzDglpT/iTHPOXoRk+5N
GXaAozVIrMnFXcN9dixbV6HvfXdyh0mcx+q1rrTXyJaSqBk9HEpGG43GBr3Q2ODYvDvEIWk4C0Da
PS1B0C+semNOIuA9/y6kyBtZMNoqgFRmDKM2YNi4ITbNvw6M1Ip71oP5VWFscnC2+/a33AHFpnDL
UEZL3HU7XhrpA+fJbfhsuRtrd5fSMeuOJWfo1LFCjlycGjSISXKgdJ6/RLHVrw9g7/bld5bq7s0G
fyrGiCPvxYbfyytYM0bNVToAZG6La+IbLlE9QERC+wiPigt+LPz2X2bkySd0GClZaF9sidshom/q
YEd2BGZVuUTFvpCts2dSPZoOKwCNk5KNXAG1SbqbuxQs+WZiXY8dCzghaLcOIur60ieCnWqZ6h+0
obu+ML8F1qhmhasOlBBMVfTAWXUUN5p5Ht0Ig721kQaLf/9EUc2/7axY9XcJcDWocC5p0i+fjmX3
XSc5bcrzqmQlNYnCAlr8i7dRD7u5vAdPqtmm/lxhF+BoMjCTUduymxjXVSHBqMn494/T8ABnS4w+
HbQexZd+YyJqnwOjGgcK9c19Yndsk28rQnJO31plWqhgK0CggIsJlAtq8ZBXqXT1+49SQVJEU8M8
CpCGPH82vQX/zN/sLNZav68+gkFcusGdUGKnqANDVKMc/iTezrUenJkaGMpVxw7g58IOCsMQerbF
JkQ/9MQIyfzrR7YSIi5QnobCIjJYaKR5Thx8al+yuHDYZWyt1stS7Ml43hJrbCjAMY/e0kAVgBCo
YdXBoVYeK0TFZY1OQH/cB89mu3DOO9F+/TO2AhQ5Ug+M8DwFRyXtohGVLceSQ5U5spyMLwmIlaTg
z2CNAuT7vXkqr8OKKVzDnmVagAzZETG2/byLj9F1ePgLjIHimUBL+FDyQYv0ZxHS77GKpTvRDAj2
JyHRE8SX1+N/Pih2kZz9+3l9saUtqmwKPkL9m1E2aTjdrDA+ARUWeJ9ADUokalxgt4PZgAnnLSCW
Om0EKA7Kas36hWRYb0YmsiYWUuzAZsnHzMwEzjFpHzU72u+H/B75UDtRNgpLnW4UdfBGi46nANuS
kDF+6GMpQX383p89pYU0OmoZNAR/f944p/KK5iM91jK8DRSY1L4ZwhjuTTxw25TrZhYIwl7lDTAX
f3PVgEGjYu7Nz7/nEOARk849B6x/CWjZ+oKV7wAd7Jr2NzeHd+mpY0J8AHYzhNGYe9U2bBxGWd8p
d5i0LjJbE3+mazVAMucerJc6tpsD0EGaHGPt1n79FnTieqocUY3UMfYktarBLVTCLFd40AwjQTx0
mYbSXGGldJPCJJS/yvUBFZgdsxkb/UA8OwavnFsTZ6BJtmUcHaM+qHSNqVDSkmG0Z+EcS2dRu2QN
3zqJVAue7WPKgVGiC18F6VhUtWtTHHv6ZQzNf4Oc/bhvKA2p65cxDN38yfVXjHZrS/WlEH8xWIGX
w/K/SKg9Z3fIr4JJeJlliOHUgyzmZo5vvO4m3h4rVegDklEmIs1STN4meb4LhTCa2WUMpU2FFuyJ
1R262QZ2r3Iyj2ENDHl3GN3U4q25slCANM4zaCraQ3jj7wVdpbv+J5Gy3IIGz5O8+85Q467eaJPm
O2/3vd1knViA+nNTgd5UnHNt42CkWZIpi29BY16OGtySLnxRzexm60y+hxkk/xgHLzgeQwlgcNAg
5T7yhofQasq64erNLx27BOJeAkTT5E6/MaSen42Bsy5ymxAC3+bTNMW2OJ+F80hix02gdk/b69d4
aYQ1cOQO9XdYGd+iS4hrjC4Y85hrSqod3O/c6qGBIxuvAP8LWwu7s4P40uSM2cR+w/Oc1p0k/iEu
f3iQk12WCF1MvsiccVGPj1t8ZZvUW2+UzMULBSyRT29JUtiUSK1VNuLTGHRvN/3gIA2oM6RkPvnD
aF/TfSzSNdBeZXJhNoc0sH5pdA+q6/LidxwwQO6IQMJ6eeMLF2EdEXkJGG/ZJdzM7gfx/AHcjgg0
OUzNJE6fgDpAeaX0xUz8p01dXWIiTGOq3CUGIXVKJxPBys4rn9jlhAMm6EjyOc7ZoCtY8ztAtnvU
cblJM+kXRfv++DgNptyNyIeWoVNEZKpasNtjci1XBZMX6k0iubQwwRpTyqsQrRVu3EV9XXdOMm9T
iHPT/i0jE/Lao99TIyQPi75LiGu72WtsP88fsPYl7I9xz3qtvswJhvenNzg0lcKQe4okExiqVpRB
a0jL1zXn6PSzVLmNJH2H7ct3OiB+P2VWvJGqkU5ul+mOeImT0AvQscnLzRWnZiRjdIWJhBD92CRy
tedle4THjke96/Jx5i6BHaQP90DIiIGKTRrpyoi8pgWA323ZQIFtEDYNIWjqiT76eme/gBVM6ho+
91DMKYAsBgiPQ16hEJbWXS3S9YKlX26P4fLB3MyPFCy+Igc4C7mGMo8ekeGgAAKSoEI8V9Wx2Zps
Jxf9e5cSMkor+1kP2TPdmpI8KrvKmNXeCSRldEC6V1KgoELL6zpSjOqR2/FSSj90y/xwE3AHWGPy
zxFXAiNx93Gxn82qBLLTFxDtAzdKtk6Yit5dnHKN9DAF1EOgyBRVTmzR3tSR825bn8nWiLA+wFf/
73dBCvMelh/Kk/hGuP0DuOHpfxgyTmDycCBR4t5A4m7lXd+FcCix9Pt7QssFJc4VGFGL8oN41SQD
+y/mt953UEpmY70DdqCCt3aSo7edL8h5pLCKRSBKmc2ooV5bKAxJOgZ5/UYbpkFI9pcK7N4h6jKJ
K/Doao+6Jx82L9r2EZb46+yRSx3W8VNsjgA2CKR4x5LCgzSu1RNWLSl0FzMt40KWihdLQnOzxHE8
EedRveuhot8j48scVyhGRCdvtu7RYXUxLxroh/z7fwFF76wxJME9eG6w+nprIzZ1csziKc1byraV
y1FZKWRz0qMkdTs6em723O6qJdBD1p7pxi8YQLcsEE/5w80EL2SDWEzCy56NwJbgt1XeSxF9cNeQ
v6skrvyxNSlmfgOms80c7Bs40cJbr41jIj6M/aIHHd64pxacJWszcXUigib8qJeVK+ltSHMnQjL0
3MFvpbPwIU+bNEN4JBzB2M/tzwkc1TRGC+6o+64gez9wtAFOPCOeU20dCfdHGGyGVl5Em4aU+LwY
W72cOjr7YgcduoKiX91sVYqgguwi15V7m2LAinXzdHOnTap3uNQ3Y4x/kTwffPACKzxplOV4iJBh
J6zMRu4j5ZHj7Bq7gQ3MQoCJgqjh11b0PayUTRC/JlsFYAcToOsw2wciIznWhi3iaodYSDnIuNey
+dvkQMNv4jl72vaGgIFebttMZOl/8yubYUOKsbBmvhSi7QKd+Ic4KKecNxNPvow+CXUISMcxqTGa
86GBX1W+rBdxt2gt5amaG+9ZpsZL7B1wDWEdyDoOajHLbEBRQ6eBdtKFXRWamyEwKkCfXKqIDwoV
ndlml7neQjwSzbT7D8A7FqJQDgJjI5pn4ga8TR2sjVkddc9EbezF0HXFJ6Wa1P0yULzDbs4YOIui
9VMmyuuNSe3J8sH0cQ6KZblytrz0VWVBhY6cDIbXBxz0K281dqxM6hwZwxfEzW+Jaai0G1IsIsLn
ynV2WgMT/HNXuyLbiGBncYGPPMEGCj5ovM6x+NacUHdeaA8/7mF6WM8qx71H9g0Am7gc++12UHUt
cKBqXrTLmaRdLHQXXf3ijOoXmNaKpv67tKUoAuynFNDguDG21rCahYPoclJm9vPYdWbr1aFb017f
9C3D39gguxBhuK9AAGCQkUMFIGCXNXdqz8/KmG2h+LKYTB3UIKj7beXF0ikN2dVnvs/gA63uiAlf
JIcPWXhvQI4OBP/lK8qDROycuTCrhugHV7LzC7TqPuAXMO2W8qf+ceml5Xfy8CxvfhMoHL66iukr
KNRGSo5vqTPtSUGrB0XHrvS0mGsxXnU4hcarEEF/MIeYfazpwKa25bqXMAWZa98+DCHqm7lsgABB
jEdaBxUTuVAnKifXzc4ajMlBeaIQbVHLTM7j0FQSR9QlQps5dw82mpJtondBoCSfRGg9JU1/et5U
lcWHhgmHcAQc/4fyRt6M1eHG8r5clWnmPFCiNjFC1NsZKZYCWUF0q5D+EI6Bj8qIa4cAmN+y3VQM
M9B9nmpQX1zEky0WY+mndJVqi+aH2lZT5ZWeFyLKaGqZ6HIPRAmdF0l9OeQUhJuebGQeygEWv9Fy
qJa3mkamqqj5Y/OIRNqLZfgYO81J/H7KV4EhXpPrVE7odFpya4AQK4Y34E8+9pGkm+FkKrZ0OlyQ
q8gQjcznbGqIE7zAajMeYQRMt7KOAK5QaufNW0pRwrjlEab7aj7/6NftjRUxjL57tcAgNcEALssR
ngHmiJc1TUtNmViQ5oujy5ZzyKtGf1pXOCABOmmjlLojhfm6N7wLdkkoALAOUx/r8dMLmCNPxD56
Sw4nHcFW/CSj2kjfw16+qmlZReGmf3fSCqwsiF1tVtyPvzKk1uj6/fGPKPARjdrTwyNeIHOCM8c1
UVvGte8AJg2Bn+UCiXr94JAyLTLHPnXy2Wc5Q5qldmDaKTQGXAtU2A7UrN2aLLSM7BKXmBS3gs1c
Jx7g7xB2ijjnObERg+KnVhuyIkOQV+doer3xV1jxNOJ6nSDPkBtYQAgeK1OnKd68cdRibsH1VH+1
437xgxr8GUR4EDbhDo1VBzYdgPuoHfF9SpL/b/VqpFUViPbGxoYXgeduXH4EYqJ/HMbCjrF6JO9z
tBysClkxE7JnnodYB33MzkdqCm9N6I/zgIjcBYh3w9BUtlGnlZSGgeCudqCM0oDXrxzvogE0odfb
vAx8eG5qryT1L5CPbsayPzBjVUR2TIQz90TwaJNiPyQUtoER8LGamfDGm5na2WcStPi8sv1e8928
h2kK2mXV3bOVkGxVoMgeo2hc83C2kojn7UQQsmMzySeXZNS/5M1LZSJZkpYe7QEmwYTvbohqdONv
sIHwpQk4N54AHd+RYR5fAbk2RL9+cDAWk8nPoHJPHYZdffVlcrD0apAs5oEQgAH0VNf1vClKrtaT
896fgBvB5/Cfdus1msMHtNIbkw+jr+/Y8bloE6hmu37tacHsMRQEAGa8hBECV1f6CLa3nvHRGL1L
2PXmksPf0jAvKiW3ODkdyPjES2XCEbOb1c4d9/ad/w4AuwrreKbKCUtkzM0KVpgCVtnroCgm89K1
2RWH9yiI1e0kSXW0LqdQWNMvUXgymTprvC6onQaIKKVzK3K2qEwcwOo/YwB80zXkyn8em9PIAUF4
Bmxa7ABFnj1c5Mc9VWlDtDfIRloB3FaClJX22jPLrkMVljxLxljv2HvxsJ01Egb+0Asgt35oufKN
/6gMa9hH/4AQNCputiUHa91nrGTa87J4r8dusPulPYQ88tA/eQacnd3k49ifoLXrMIBaTjkd4IWz
gL0t4ny4JaOwls8jsvJIxTSxClHj/bhYT21peRF53BRi0E67V3m/s9pV2LX1ONFzl5yIjyYxBYTP
WfAAESrjIEsO+vTkOTWfGBEJTkhfIh2VodmsxDqYgKtaEnbwRvHEFdjWjS1PNnygUMkWWxcQLvr6
Qv7OTOxMgmicmZFOloS/eVyoIdaBj8WKnE11UBHS9UHr9I6+kDN8Da3BhqCmJ2HsrirA6hmJzC+9
2yhdKaA3+CJI9Y2qDu7gtlIxCdg7Izow0hD3cAv7wcurOU0QRI17f1sur7/XW3wMtUGzvQ1m/c8B
vr4QHDsDzM6oZ4dT7CIeGll0qaw42Tpb1evl4zRDPmBa7sUPegYFc2QUp/8n8zpYwqAbdH3voLxR
aEwkFyo8RO2QaKJU3nVbjr6NF7TrDpaqXHWjz/4p/UE4+XRNnO0HmyNQTp1Rd+VIv8UAFyUKemZI
afensFueN4XrLfDslFbhZeU4jRb0rlL4FWcuc77Jq0TjXyp62vZGRUezCAcU7sjS0z27OXwzEmqY
XiUGeu1TIMif16qdjVyystemWF3t7hXv2fnvgkgDsh2toYHXPpWV1crfA9RhDgmTn2nIY7A9SYeK
FeXR2kJv9p83jRcIdXAVJimtE4CDrAIPnRP+zMkhabRHtw5GcWvmjLGRd4HpAjQzb6juecpDiLOZ
LTn9EKp3uAj9fqO5hgd9+Ywc+YXULG0QKFvxzHZLMiZ5zTgNnMT6XRaIbdUHYlyQoBNaB6wzW4mL
ybOMej8bW89f6zjhKdYO63za17fa2uozOCQMoGBpw6qPpr35CH22UEbjOmYRrd5G8lZTI53OIsr6
IcvadyIJyGts5iAsyfD+sWl7caxZJvYpVTFi97FUsy02maMD9q78k8ORX4ZheNmrLFvWdZvhD9bI
D7BpYyw+f/8fW71zWZh8CNbVd867L35kUIhaffuqXA98f8iAuD0l7HxJZjO1+i630LbWc+jJdnM2
GnTJY88NbASVwizZe7Jy7Md98cCFxfJdqBgyDqe3bhXxjseFs/4lqSLd9a0Pd4Ya7rv8OMNDs7Xe
BHOW2W0gPDtMmUAjpmLxo/BIGEUDpNV2KAGaKvag/Bfp3pXRGXrEHY3iZ97irOK4cYjNhPLuXPpG
Bl+tJJJvHbCz/BINloyY6UnUdOcYN5dz3zb7rnM2iYo8y+H29+K5bImxHKv9tNs/wRFcjbaCSh2J
RVwoVvhR/yzQARlvmRplNL83H3TgEThAMHXPH1/XUVpcYVUtW6kAf51FnzGz+wh9PVn6gNilgcYF
z5lsELa8CnbVjksgkq/5L/3DbFzRqTS6n2jeqaiKudmOb2/G8baFMEplj2TImeBki7HPYRmqF5ji
6fPtjXT/CABny/WfcQ9RUwUiG2nkZdFHAuLzx4UJhgQvrLNQH2PBneZMORssZ8d1uQTIgTpcFJBm
wxwx31S+QIu0WI/ZI7SCm12+g4Je8ALULwfkugP7T0HfkH2IbX+h01x7LHBiiqRc0W8sRre1QPDs
ex5a51h/hFbwGffts4Z397unxCKy+nn6vNZ7dXx+IbH92tjNsAqQRT7o2H9n7lGNfO0N3Y/L6otC
hBIbd3qpkAhJwqVj+k/8o0TSc29Cz1zLadWruBjwD0tqV2QFIPc74hniSqx6u0Yymd4mLrvpIplF
L+eTMcY5IKDBeRJzC+gFa+zwZPp/OFb4aQ5t6VygtuPhR2K/tVNe/OcGXP2gShEuLzpu7pML7gZw
/OuZ7zyL0EkRrcGmTVrgro1qGliYUd90Ws+spqT0VQqO9XMApHNSYGsu9JENNwqYNvzoAGUfLeUz
pfAsKoQcIL59sfs2Bz8XkKnMpx112t595DcEYrJxlIRf1LlAq+8SuoQZyyty7DJ3vs7rPsC0w9rL
wFu0YrE1FW1H71xSJAaM9rNxH3P9ijAXZQXb9qSktEuEfZd/b7lMJ8K5klB4WBlI4NjuU3KjO3JL
5h0hRIzgSIn/b5D84XOQ2Zs91ufir5bOgQVDME2pLqjwzwIf7TEdnanl57BVyqYjyN0qqdil3ga2
ZSkd5WmN5J8X1ZYJKFB0evFPnvH3dLCX53O6c3ibby+rzuUPOYX403ty9PJfqPzZTHbstBjXhSJH
junFV3ycAsXmq5+ENrOA39shdCFO/q2/P7JsDs/R/QZ8vCZtiEyiqT5nLpWvQ3YyDd68+Mll1Wao
TBHxN0NatnJ43HPC31aemjNH7r6QFJ7gpb/6F+gH2k/2/g/+Z97W30QlGsHrvlIPEpC/d9J4HG/X
qfjhQ1tQjGFL40stQkLYSiIFaPkBvIECf6gsGJroe9ElF9IbYcqQ6HiAzvzQBD9BTnTzbZHcFMty
EdDDG0vXf520nJkwdWifQnt3SOr6ioGnn6etqCneJoq6xuj+liZP0MdAgeq34KSuHa3EshcI203z
D4mVvjGUWrQoBKSWTksVyezJUEtvTUcTMJnBDon/KImK/ivvUfoncQpFXHO5RWb+Y2nPGEPFRgCv
3OSkIbsAgDZpheI7fduAYBZ/xizNWnVC7nOhwDr64j18pEc6hR3IkbvMGViWswQx7oB1urtw5bqQ
Lvdhq7FgrepO/yfi51fZyx+o+15CMZ5I+c/N2aYwemxazEJnQ5QCcQpmoLqgaqYSCpewmdOvDgo8
4kpMaa9IfqwpU1CC0TLXR2Ml7pxORFi9VL0IaaMLrLbXDiMiDqelcsOddkmzT3HlqM63wySjAfUP
JWJEs+d9qMIxznxG0UX7ibD/PQxShzxNw4BcrVhSWxp+XiYotaXpb5mRPX4cmBV9NGITveg4lxeY
6RlJjmL0VqhATjurEirRWR0HNjiWEIhBJ6/fFI8nzOkh1X2ZyxdGHI4KR5VcPzgyEXkwNRrgrIaK
NQ+/sli8YGzJ3bP2+1G8AieCLQH26+Upa4jPtiBAkGlL7vCqfff87hBZgV3XJb5dWPmmL/oT61H8
gpPEoaIY3NcNyHavXKncxpSUYLtF3AGktBpZNcvxj7R+VXWGsrQNYNHJLPXnpKBZvSekJYmsQeIG
zFEl7FmOLQf9B2pop26r4tOChQKr1EFnnUK1JHP9z2hfJhN/ykn5WpIzRkpP03cHkQIFRoVEs0M3
9LtZ5/kRX2mtXbjZRu3no5scllgNKTqQy29oCE2Q+IkSZQ5xBzQBrAnSPNpekzdVB6HqcuGic0Rl
4PKUSWTUSwaeM6VMZP6iomHWMeXVUecxglHhTOc4amDZnbwFFva5h+WGEQQzrPkGbs2MVmVybiGf
bWSY59JkDFK0mdL0q9SFusg2lvGTbH/r4tx3yFUaVJaTVvUHh6UpMf4GN7XxOWYtygiQD4neXFMO
mkB8AkHYYPDMvAJdycqo6gc/GuebIySOlxnoK6deZLyhuiiViwWx5PYLyBE62wtFymIqehcXgiE3
JfQaM6DKgCvz7cM+YjsN1/QKHscP/KSnrbsi6TcZdwbj8yW6vYx8N3G6Yv3LvdLCMdkU3379ppgL
0hGwzLqfyVWfF8KoaoBUrpwWkbJGevd609vN/sCTpdKmmT4fVyW3rsSewm3F0PE+NG/i7d1JiAkk
cqfJeEMS9bZJJwxCTsXQ4/l+Cz4WjGiMBa/FkWzPilmPVzKOw2N+jzia/fbpcPoEJS9QZtpooa3u
3BVtpMqsV1NlHmrxKnhjAEisJm1GHC6rRZbhiNrYjoFsHg0Wahjlrw+tTYKkq5sEGuT78WipCOd9
ZL8DflziVOzLSXMu0sOdwgT/yyt3OTzxHZGHU/DtzBmAf8nmJfYJ2Zg/dfYgJe3TCQYDeqrHBhN8
32StIxIOPomvzluJ0Izn8X3t0U7JHdPd168tDIFj5K0mX+OPN2fRRwLSDHEWqStxVLlLgDqbOZxX
g1Rz+SaZ6B85UShwdmJBEYX4ROgxemW/b5ET3oIQDSVoFit4e08zgeGsdzhqCJhNFraKzgQ0lP/y
ZbZdmHsc42TvZMx6rZw7g6tvE673A/pjb+MWO+PEnC0adGlIVIvAus1Lqg0H/aN4datv7PhNSTTz
d40+y+PZdVVFY9BEKybKZ6fxdt6cQXNt8IxAUschX800IElm3GeNhgFPAPao6WNCZpDvJEOEJmlv
+RVjDZw5Spgr8RzHcZnF5Gvs4B66wQVLybZfyuf59Nmngria+E28u1cxQnYIQONB+N5BEe5Ai+35
HfDmwK04HFOmJ6yosBT24ZX0eVjOUDsZfiLinYLOOKmCxKgXvThZtq/rGynzJAzHyP+veoYowyqj
uqzMq+LBdBdHLV3fhSq4cn8/tngVg5yqe2Y3k2LYopbnJSG+yWrZzatkjqUwgriKbeN/A3FjqAem
vqIU6hfzubcjf3dL3g2xsR6pE0Z4t7UXYtU87mYvlC70RoSHUwJ6YN9s2vyTQRyWo+aty1i7+/Qx
k7wl6PzHZeDBrZ3RPnqxWUtK4ZhVIfBwbEv4fhklItOJHvqMrtsu22id3qv0XiFECXdZJRMA3f8S
MlDmddG1iuhH+yrpmfnF9Htt1wLWi2rLWDFj8fnDPJZ+BiIGxE0vs98imSKTgbbgv+tnOzLdSjc/
eM2dgMCI5GVs5ld0pU7fia8A/MnxHJCU5r+J3Mc7SW+GEtnNcdCMADs68/vFBu/qEe0PuAoipCAM
cbFq+wtQrmMA9cZQ9YqwkPOINcCfGRyVn1YH10mxsIEqkZPplsyaITwOvbGv0RlsTZNnbk8DVqjF
dwoNHoWBNWYqDZaCustct7dMbqWLWC8AbPBE2Pbc8csepm1WA+U50M3Jahiim0BpUuuSvaRzcMN4
Xw8LVLP0HJ2jYB3UjYoA8ZdBGO2HeD/zVidEKw5y1Nyea6FbRy/FcYzSm5ZYSvHN/SKAEdUyNjxL
WP50MYUwkmUhAw38QiS76FP4tIi86RjrI89FHyWvnyTPtEc7AH/TDnK6VGXHQ8+cma5b1mdSmP45
wg7+JQz6PH45lgdS2Ibp1dQH1GW29tpHeZwtj79NTjTN17rfbIC+1ULnW4av7/mKzEJmGM1beyvY
P34cchTuCT71OIE+AR5y22ylU8CJsqFXBDjGxuMuMQT46xUC2b8x2U09qRGR8U/8JbTMMuRaZGa8
31ztKOPumJ1/cvI1JbUj+3oQrcjK3OJWPz8jGzsRgo/9gBxOI3FEN7oGSjP4g46NYc1ksVQCVaVl
DAnVpgLCALw2I3ZRR2frp+6yNwxup7Q/r7nROY/EzJOE1K6lEhakjNL5R7gF2mQg8G3rA7CaOAZI
C4Ntqn9buD1v0rGul4Dr9rDfSXwPjQSwJv3obZM/PpI1zWk/G7DoKvHQrpXOTNiqDIjuKA0Y3hrg
qRmN/3xw7V4BayyL6lPPC96knsJCSwWrGFSVjY/QI59q516pT5EiXqPNYJhTP/zkODFqvDhcsvDq
LQM/FeSQI3tmGUjO05SESbyFTdp9nvxL+WM6uhD/3Skt3XXgXeoaVKTRcbOJO7+ehmt4ZdAa4w/Y
H0dix2HajmoDSNyKFL1twLE4JJ2BtfjRyssnVIDKrICBx9B3+HuUjl0HDllUzsSmeoZFnrW/2JG8
lTk3PH/m0CFkSmiF++56cojf4m9TtK2RJlTitJnIcSFLTkN+h7RLteXM11K6wccOS8a9ATQEmLSF
oN/YSuIz/DDi67k8NK/Esp368bVDqXYk/6x1JFqYT0iVzWkwSaXqimtl66xpxCBmN6C+OpZDXWSx
l1KdjgBmFtIUclQgXoBbItk+r2hMo/WqZsQ85BP/i0HKfH4KLTqIvP596dZRmENJJO2ZneLJG7vy
tZx4ChCthjTeNiLf05W2b/yKcaGPqdj7nNQOVz3Z+PGtgkCt7zoXG59Mj9eOCs46delwqSTsZE2j
5b16E7ZKhUVefpbh2QHtz+yy/UYiAMQLIz5eWzK2sjmyLuj6uTR9dDpsl9WEwie4FWPFTJr+/d1o
Z705/KIo6jyLVTP+bWXdO8+8NaLJSNC+EPkhPw7G+4EUjsRGXnZDG8qJ64aKfWtYBhhkvnlLMHkf
+AtL3lWWlbXdBYCykrKlnleg8cqaI9BoVHKsSWNJDgIkXyhlCcI/puOdZcaNsT6nX1QImNtu/iQt
lEWlpsLYH2gL1agPkGcn0x7Nn6iXJBRX3EedIbrN3GHw2JVkZBcJS+ZsRD/13PF6dBwGsZgXWeFH
k/ZXf16B16Ob0EdIoIiKO9NNj11NQIcpMQr57tckEAurryczvSe4Dn1WUluAzmVPd50yHbij62Cw
hSKdU0exSSh0DFv9buMgPXO7dYgyvKWq/9b11bau7OPZkWkknxI6KREE3Ufg3sidMwIgllhF49Or
WCGuXmgQipsX6CqHGxh0nLq8RUT4Qe+yIcF1bQBVtQiMpR2A6B0YInOJIEb2pIByFowyuU+UVyji
sw5+sEOJtVnC2evtQj5mYZ2BpfRo2QI2czK6LXpCxD1GSuMyRceh8DVRpHRBfYuWHaeGNi/dBBVh
zPkzTz58MW6gAt1yuUAVJbyp0zPaFMpkQ9+HDgLRbc2DjhecKpLeZ7ftA0O5R+9Ro9q+Bbkc+dKH
4KH9uSuoVckqe8SZLKUexcmXSpFqfBWKqWCvcocU5aMwyATeIW/60mcL1kIFBELW+Tl22MzP1/au
eouVAxeVQ3MN8bSyNbEJU+uqaR5h1TAYg+FsSwlf6q0OlvjWXZQFjCv3Z4qFtHgmcf1ABFDn2T2l
+DsPph+CMYAXmadxQKIo5+CvD99LIb9KpCFifLD4utiwNgsxUCP4h7vs+l0sLz/0atRhnSa9F8PL
azY6tFB/M8EkAZW+uZr9NE4fVLrPJbTzUDHM8AEQ6xdAuGpNEZjvEBwCNvQoL2fCcWz7ZAgZxWwt
Ffgbijp774EgR25EkUwhQ6DIRaAHy+NOrJZ9rMCLtJcWrcTOqMen9/0QdB8J+der/368fxYBKcph
yaTYdyLf+IkjORYljE/ItTp0O8yPG7zmG/tAGTDsTR+QFa4FML7FcgTCo9N7RIEK8Y3KESgFXt+z
DPh2x5XIZ+MHCmo1s5B7ERNlbj5Ho5T5YukUT2gWWmfGhnja04e3Jug9UVWg70jSPk0FabHQGc83
5MqZdrWbSj7nTdhoCaxUazwbdfMevinMR9UhGckfR31hWOmCZH3kdsq6vdy/usxVXCumphc7dlfn
S3L/TzrZnUXJIG6yPZRzCCFnld1naynWeu712giMubocRK9LLQwv9JefecjISBkDyjsuCCtrO7uL
xDAl4WBjSJx+5INdOLbUNNP+0vlILTMoCusFaNRYNT/lTBqv9g+vI3mn5KeB0KOo3hY4FHWM1pmS
eL6bKoAnt6M52N4gHVOOr4OM7xlrATgyPTHKCTFmFcp0qDu9e+p8t/86fZeKmPwsbXaDvj+7xxzn
Kh6jWGF1+sczLrhK0JUcLa56D7Jx82t5M9+mkzCLKbiUChXaGOhzzZR9gI2gdsDxMoFxZ96XR32E
9vhgqdIQr9m5VLy4moJ5toR97tbvP0JRuZbgCn30LNwPGE6JYLwWmSNf1WQX6wgAaytZzwFsB3jq
0nhgwdRUXtLXpkIPQnwwKaVkl2pBbVNAz4ThyugFAOqhv1pUCUTyOq0x7LQKloMJw4wWgtFf7P3F
1E98XtrClG0zcJKBr9LQ/I/9cTFsyG2Mxq9+vRGmJNkUiVmnjhjYP+Z8BSSaYv+KJL5cUORiUgJ+
wv/R0B1cOXAyEegVsvj26wDWo3BFSwviHtVCoF11mRV0sz7VMX/UHasCRt6f5LKYCdxURLaLxtzk
DeH6/Bw+U9ZIpfQkzW3Q4CdekFyXmG2b1M8GVayPrfCUtznTc2+xu7TphtWDjKeYc8CSJZmfkgrG
GwaRjO4cEIi73rHTK8nO9CJIxB5bHfvd5WXMqUOthh7iTdUC2N3ZHkAF4WAtdk6vE/41rRTllK1M
yCCMT3oyDbt/tHfSCDQXLOAMxPbgNIGY7ElaDDVICBqmdEiavTwW+OnefAc9NoYAXdYqBmZslMXq
AR3rQp0+rswO1uzV+JR0nJ7xDTspyz7tO/MgrCLFk2UHq0vKxducgAdIt0+MEiZdWPylslgcJp6x
ri/gyQL1QtmKvwxk+hazmQ3eRWkY4gSwRJmpgA+C/FB70aKIfl2URBsQNET0cEw1Etm3BquIhDtp
IOHfXxx+B0JWGQOWfSicVH10ZDM4Iyn4SJTtq/RhhtW+C9zl69dZdRzzELRX5l1B7tSUPifvD44E
5jRxsyvBnjD8HB6nf1pmbnXL20MMJZNe/nBNOzD1XUFZJDUFnCR8B5/LlMSnoZWIF9HPAEdhN6q3
soIwYM/aB7gb6FiZ0mprRZQiqvmDipPdFYg9FY3jOovjwWJmMYnV+uLDiPkxeBi2GXtMt2xDfo2a
ONXundU1/kU6W4i30HLgxifxTFADU1W/TaFyWc08eH9bt4JiMjTcVq3NlgLuQkTsBQKk/wla/TVh
T9jpT/rQD55NdRt/fkkBW+iEiXjhr9cBevUgU62swbhS5zWWhcIndR8rsfWdCAM+ShTFeH/xJ6H2
rVFJZ3E3Pq1DTogJHpiERZqP5D/ALRhu4IK0zNYP0rTzPs14rOCzXjLSHRA41Na/vrLbLjVaBqLh
7ZTNbezbcDk9hizKAsXKShysV8mDhM5+tsI3dwftRvpgabJGQbqkhSJlnq95++R8JFoWyOjCIxTK
zQj0Cc/1hDseFhR6QunR4Ph/7W30w9mZM86Ze/wXPWEgPF2k0sR020VOvNvKPIAXgk9X/qCPloA9
a/wrM5FgxtuhRsu05Lk6nJ87nXmAfIUUyqTYgP8XV3DnOzXuaMhBOeXTUt4EAY9hm7xk21bVmDGl
6L8hDvu9Kmc4s4aCjYRAJw+FKJFNNYszWOvGMhmwTBvhkOBgfcdWn3Al+bRIhJl0jtOG8e6MLIkk
8It5UhpytAGW+o2cNpwhAAfEiHg5X/mzDWOVbmtPMwEZikSv6MEUKqVhQ825wriFUE7Le0Cez08k
hLbwguZpEZM6pV7w2NR51oP3GRC36HSZOy7lnxGM22mZSBHyD1keQP//48SS7xz1Tfo6B0OodUIx
br7QaC6DsjJI5O5SZRZD/FWMpP+gBUfqMalXUyabtaWJxg9vatZHemQKRv9deqgoAsfue3+UrMk/
0GWjZ74NIn+g3PMvh9lWRfilkLs0q4PmnquQpngFL/kZBegdiDu4urSEEWqivCBoYGp6SCC4isHF
T/zM6yuAKfxXHQLm1vSWctWUNOsP+fIWF1p7cRvUJq94Qc5vSE4hapCzSQBhrLF+h/CSmBQD4NOs
AnRKSGTOUcahbcwWLI8u+AcVjIAO/S6lgGA5RWgTdlVz5TZqD3oon35xEhZSG2ReFMTfEE0fD/42
g41VswooOy5NzfkTEYLyNrZU1wQKFX7bqnE2vf0Fd6uMn4mM/fcwhoowwE3y/aZb1XRNrsbNmOf2
8CMvGK+rZuzog1IRBaFuoBuCAPpKOg6gctoUJzC6AaOhxoq5UWmeWQ91EJheuIA4byJZp0ldEy3r
fzq15JKTkDCrL41qrA5FpHSVvZu3yh83B1yDftoSaqKYzfWU3x0HbW9KRqzHuxbvjFcnXgDl4mPc
zQ/R61TC6drpUkLidFVpyEvOW9usMPNdUbXELabWhBbWNq6gX7O3FS2S12I41ZrbUBfCAf6y6+ZB
fWSjdatARRFrckEbl/lCxtS8tCXTsRSgci2HKQvQDIb8/OQOoBlVnsCztJRDDy6I0h9uKHBpJL9i
swPlSfPA2xSTLgTavmdpmyL4e4in8kkaGjfDwqmswz+5n+KDx+SEG+zreF2B4VxbiylxajPqYNU+
sh9qURbnaJymrbBCPfpgoNtZFgX355pwrXpT9/ZCigHJOwAYtIQZlx7gqsfEULued2fhZnPjL7sa
IYx0m669XdNj/s52Shttxu61B36G/wW6VZ1/7pw+YENCwZnNmxaPJ5k8BZnHu4mANhWhsP5v7Sa8
NGCAKR4F3yZ3jdTSKA5bvjBIbCLGW/lWfBAyJ/4cIqadopONZRW9nS9I76S6cNBx2OlndhqkONBG
8hoB0U1jCCi2LkMLB6NDzo1PKqid/iLy9q47iWdCM3k+A3x+SjztU/fnr6QjB1ZAhOsolb27JOpg
yBZZn09u6h4AcA/ngPm/i2bCcm5QCYtNxW7TSGrc60Un1KdyaFotxoKxbHaABQ6P3244H/cAQtWa
WJXF+SZiV72CjXlBYUwzrnV1koZpQ7CTbcUEXV5a8YN2Fdd4+/c4TlA579vAY2W6INxIGIPELC8u
G2jVyF5nlgmUUtEKIKFUflVm8TdgMW6mAScvvCbbT0xh8E1advRuXRQSEKRHN6Felzi/6Dj66YxP
iZwEbOdCEC+U5YCduokU7RTX6nmjtaj9nASXkYlFCmp+dhZYqCOpqI3i4PvXiZd5VlWKgNSRTU6S
mBLgQb2gcRe3eTdrmz5RCvcJmMGsCpD1WBZObhPODRZtQW4/uox5K+xvSCPuczMTY/vBhUbU5tbX
E3Mo9dBvHDxGP/X996tvtNQdblPb/gQp9TnHfuU9wpouWh5nOKkr/faK3tiylpG6R2xb9l35XFz8
weLAvGzcowZ2wagW9sv8pqjDaBKzVZhRXYoZndvzjV2NKHAy0NTA9iKqqr5hmWYPr7HmCr59nygM
BNQshrL1OnfvgL4JaujpIDB1ENpu9xbz5qnvukJgzk66AIht1FWDdVUBuOwtjqp8OVRTsZyrJZqu
J7yQwyzMnDeWC78zTT75Srr/GqJWR++aX1/ewkvmLYepMkat6u2bAD9DI53DhEwxLIxW7eIXg1AN
057x/iLQfbvIuYsEASmghS14opjiaw0d6O9l2R22Qhex7IZjQpKYuvF+Rg2+dM0GjIxrSMC+lnEc
TAh8wK7q9roPx5iDRiSx6ERifzzZ9rjDvEbjqs+8LrgRbZyZCTL5h13hD3zbW+VtpOj7bQ3D7Ppz
S02q27czyzQ2JVrqiVcl749w/srOn7i0rGQCsznwW7atmkDXUrSQSft/Mym0MK01tE1vd35gc3my
YGKHx+nRVE3GXYPlNTv+JIkUobOKSzaS0yk3i5kWvw5rh94RieJVLfCI0R2NsL1r6Dy6OsTVPAFV
Ezd+fy8r6Uv8iLMuwP4edXaUU/AvTz4tc5g844emHXqLwvCs6RGbGvCjHCZyvmsZJC20uu0RRcos
2wv5Y8YYl21/tmSTWWc5xyp44Zc0YvRWlgzVd6/+voaUUDYF4lhbJHKsfT4xmaqGtNDDoDpEzE7r
mmhDewO/IcXIbRxAdmS+Ibht6SPTL7xVvqcLAUx5m+NJHXRciXVesRMqguexTnNzeY48l7VlZAT5
iC3KdYSwbx+1YjUXBkPX2UpvvcNO+1XORUAsfhBSZAlYyrVyiPzcar/vw6B//JdM0iMYf9im4c9+
KC+jAt2cN8ra++HagCwZoy6s/BOwdrWJk1BlX6ShHb3Zt01pfMA2AiLosUNDe1UwC5waaww7ByjC
Qznbt7p6yA1jlN2AuC2pi6+rt7tAmWDT30IJagOZT+c57wAroxdChqT8oYT0sDO1tNNwCcIA1UIc
YdJjvxiSDQIB1vwonPfYc+M942w5QFd+le6FkG0QCzqvbj4mde192jHU38LVNMJm2vMkl9+PKaxV
RSYsBSC0IEBIIxr9c3rJ1CBtZrzE7sEBK6buFZJJD7quq1/5SBCf9uCmswxXd0D4CXLkjuOGOM4U
U/hz2GHDr/z1gem1+idB2XCSGykxYu72fm+BigB8Ycu3gexIWTb1t31Zi+YQOgyKeczLsCw4T/ZN
gpc+Facgxq8IwiOT5KK23Ys5EP0JW9/vjwdP0TKiqcXWk2SQgg1o7gJbOCZO1pgeGKFFjG0S9gMT
3bopfN0l3hKT6bzzw5yo/G3flCBQ9ABb56YdgamLGGvD2robL98TjFTgCH/3v5NyrXhmZf+rDXaQ
eSt+AWLnUNwTcBmO4jUescknG8QE94RVFwUyj7btoFU+aluBYUY+gGuZXYda2JgEykzX3FNrziWB
JXEFHtDKlFpNxfdCcbU52Q/EEBUd53rODiAmUtXSs86YEDYBSRi2vmwNZjiVAwAqOrOwrFnIKI/V
+3XyiOAWPa5uyRoq6xiz40MHStnO+Mks5GiLBhi2GNzIrfV0ehjyT/s/KwKE3jia2TGgDPVgaDqV
JmNUiHwA49AiLl+FaXyoGStFeSRWBKnsjZqK2VTAU2NbOU+Jd5wcxMKQVT9fTRb7hhCeFAnVr+Wj
TOuB1CKrWMnEDizjhlD75DlYgDA21yNIRLF1i74H3Eml3RBcyigJvVnTaTlyNux6B/zyzkBiiOIo
mh3nlvyj7lKZtf3rL3MXUhkK4neswF6Lxb3N2lIr+k4CvKNGVPGUvUJW0Mcj4v5zLEOKR7oOrunC
/PUICDLcC4f4VWArTCaWAwEZupbEr49K+dtB0xdUk45hGlkUeQ5CaEq4Zxzpwablh6vE3SE/ntQT
o8+L3Pp4QTyEQ7qLYN9mP6wCjBTmM1TRqMXzs+cxSlR8mpdX7069KkOyQNKei9ztLvpAyFjVV+bX
iuDRpF+efwENbXBtjcHOA5UMsBQfI4oOqmr1yPJ1th9Npff9ey4AWY4fk/YqEpq5x2ULtaW4jqlh
RZLwORQUqhFrtM3AaNiAKpOZdWa+AZ3qitbiyAmE9ikUEyJ2hY3oK9mGeEE0Kk/owyvlPjHgtWie
zC56VTrNsMBVqvfniwDjxrHLYcqOltUt5Cs3kdI0aPdhH5HYNR9VKUf0Kx88WwX3GqMhYFUfM/JY
/CVDVjdmK0xYfbfLDN/6GwXaaGl5VVPH41R+AY+O1CiFsgvz2itZaw0v4himo2tjtIoR5Z9TPeJ5
OWuQd7+YB6tm3fOBAeVqIrlEZsdt1TARrYmn2oVaERvM6cFgiwVKtQ4/UwqSMuqYh6UPAtpBtH6P
YaPQXcV/GaIQMqCvxbu1a66BfNTo+vAsJoSSAGtAVIMRlz9/wTFiePQI7rCUcKwTpEy4FxBWx8NE
6zAjGdNk7Q5xKmKYcysxri/gNMnnWZiO+RDGv1AK3MolAfs8tqLVntdBStF7gG/AODhAj4xkReyV
eCY97YlWAope8qCUgfczuBywAvGGQwkOmcPR3bPXEHFLe/H9sT6FOi7wP+X1sOSVbYp4Obez29vP
uSOmu9r72ExwDrbRvC1GYAI8qITh8pjNoVVNeF7lchAcDulW77hQfYWO9X1gwLk1V3X1mZa3Weyo
+Du3kvV+4ur8G+nw/kHw9eQW7UZ3u0T8b0gzx9pwGvphdEcK7wijFLOe/zeGIUfwhJdol/JdSJrf
SV+RGEqC5poTriECspjBVosMsUM9X4LqP+wyIIwHT0FtZchnnm6RUShDaM1dVA1Wjlxp1ebwKnWe
5PlnWt/SP3fn4nCQsjeqSAJ/tSC2dGdPhMkF3lm1IuyMZBWjrh5ka3rMFab0YO2cBsCnlYSkF2jp
U8r4udnj7yd6lnArXoleRUMgseGB2myu0UwrpEUqsLjOYFITVLfbrIF1MsqNBNqwz+/n+bCm3//D
p5l12xCerFmGqVnBckSbZlMHjAXY/6fUGHopwAsA2EvmFhJ4JI8/OUhoQwp97ZjO9b+tA9+vVg/Z
UjDcFlqcqpxcsdj1b/tQkI6+w5iWsW26K/x7RqtW1QxZ89WilEL/TCvaXs3VkkbSni+/dYFZw7Fe
lXKQ5e5YtVhv79kJuHOLDqOc9BLhiJ3XyUKjGuZmRJFiFmKB7xYkD5hcGbh93P35XhW7ae21YVAS
kA2AynXC15Dt6KrChCiYzDXZ6pRKT8mYb5GVob8HISwri4mx99MRAWfOtAiSp1O2RzKFJUHgNbYT
s/NPMgQRATlkaTkKi+/SpHsoFSXOj9+u+WG5GhvMGicAJ6NiIthcejmuJyHHnuxEmfbu5rxMyiS7
YTeHzpvSeeGR6ngEdb6j0sGzij6zleuWR+JaOKmkhvKBWWY6PopEEweaOBu9RxoLlu/ihutlW4dM
xFzI8UR1V0SrF+wqFH1IDyU0uA9fItNMYyTmwnUdCel4QZzqwkrimC/FyeEia8zlGhHXzEeS5IsN
02101p8NMetGunMwblzqr5frTAtMQRDYjKI7SidJWNnvYLBf0ZXgrVg3L6fJyjCSldOC7tsVfKTB
CY9xghzxspVYquG/DrxQwGVxVzjiEwsuPVyIG34uYz0bKYHVKyQocFh1yVpAb+AJsQQJiL4vcL5j
qwtitYBq49JSd1y/0HjNFdgh472gu8PGn53kic8g4qK7UEY1dR6EaVxBf72vlJ8SF3ZMnFzoee0e
ySwcNCP5yFNuNCo/daKbAIbJr7tJ3Pmqjwfuy6Z8nsWRETo9Yxecu76nCTY7ZT8wbh6xKAep2g3x
1HkCZQYpJB4Bt5fwtPxjk8EEw0Dxf3FxOO0Pu+v4lj8MyDTWf5xvWvybrqnsRbjJbN+mNui4fzq3
PcX3sIziNLd6aGD7hsjsZyd0R8DxvbsV1n9wJcQ/MYSrkCyrswLFFxyhblYmXtp+78ROFIEVEQlU
5xQsR6NHqm5UjzfjYyDMYk57rLzTasaHwa3drndNgNTaRnQYykpMMtGMRKlPdLngK06Jyn3T/9rX
PwvPqo8LD9Jxy29iUEy8bs76amQdtTEy/lv3iKNerNHVFZdKMP6D5moIuAJ4xZlQ3Hr9yPZelVr+
k+1JTq/ocJTJ5jKN1mZZbtOc/BtV3htjnGUj4jDpk6K/s48OYgSXOZxcKJ0+bq6O5a7icR+3dUfv
w+wwOXwaecKMK0awupptI0f2JhtExoqMIcCcrvYkw/6tdH/C0pjha8t6X2ruBvNBsMw/6O83LHbq
pft3z/Ouz4AOm0DMi1LcMNAdUNpYgbPeobYCsdsZSiMZ/AY4zytREaMzLMYyDgpy5AGrySe+C0cd
+fEPH1NoHFW/DVBMnjhEk4phfMUh9TESJic0Nvjj7s/OUx6/RvYQxXqstnXGfAuAlZzPqkM3AVHf
SkfzG7z0lG/g2qr27ELyPEgd8aZxqNkdr8akv1DeE6Rc/8SWbvSxhYLPzbwXzGXs/JCptDkhLNh9
8P4X1G1rNS3/YjgK5QGDAKFoexdpEZlpgEfFtzn2F9NKGrH/jL6O3dhNLbJ8SgoZIkZx0I8UoBZa
eKos0ihyJfRqZDNtjFqBzda4wBjjuQuV+Kkna2NkUOMrQ0B+6D9xzrO6t8Uac3sasaSMyDTtSLSt
W+j4K+OQVtofiTOqoieNtXiN4/QTj7nmOBVP/7I5SUx8RL+oYNVpB5Z5yxQrBCp0xNg+O0bIooyk
8hn9mMkTnSVEBUz0JGCSgvv2U18GWyrLsyGE28/bMLHRgeFheTo5JGVFi86/cTPzeWYCIDrtO84Y
Dp6nnKruVU6wwJACJDMpGQxe0V7/yh1ZcS/jHvXa6MBjMKSX24OaepxnDDxr4p42Y8XuRrllwfuL
Wz07vXDCKEyv9ydWFEA8vXi10Oj+9PchMmKfXsbPA/CvZwMT9LLyCDcGqumy/HAIXyP6I2C9pvtH
gyYACUzxipgxQp9KNvWkaRGmT9Cqd6p2/INQaVUvm2wJjljkznwpi7cfjiSPIybzqsh8O295PkF0
cc5Dy9A5HqrzqqlrCHh1EzmaNZTFyKEpf6k7S4DuGan5OHaqjYHNMq36jbK6DB6lSD3IThhzbAUL
4SG8jW/TXUAxlHO5NTMxbqgb3gCtuxWe2ty9V1IxBk8xhh8JsBbbiEZVQUgBnqQCJGUBMq1/1oyM
1DhtKONhqlAD2n4Pl0vEK/OnasF9j1OaUXMPNspbAYnIDo38H++gNZVl76b006YINwmtwavVtEdz
OSClxUT3PUwMAv3+iSMGGZ520CU6SdjWp6vt1hFxWqxgvCDFmIO0rHVPN53IWGUWOVvV3X8FUl4c
GBq1ymfpoYfNxD9qqfJMJCoiHcywTmIEDDvEXUhhVpFZ3yRfFjpNoRBPIUOa0KbKUqEn8DkD20Yi
AsY+8Pe26IS+4o0hqDcKU5eYp4FOFrFQWx5qhXMojB715GMupnkOmlHRL90dRClwQJ1dFGpcze4T
+5Hit62SofbKzGiY/fvoeDiTJHBn45Nt7b06GC/+aAIWViRje7ffovCPlUAUgnuE/p7h9IUP0OEy
K/O7SaEenuiWgkze3dk+UfKm/EZwKssuijnd1Ru3nEV5wkOnW7ax4ogHhl0igNtuwCSMn83OsTrb
NQiY7wOBFHJ0hg45+P4xyL2roaBdsueG/okTRsR/Y4YXZ96V0+4ok0fuszMzIKFsFkqC2JFjLcgv
lwrkgqMQgfIv8h9Z56AveVzn1kgEuigJcUyCBZCBsjOhisY+brlBikitcd3DJn8E44DYT9zZ6mGI
Atwl9NcJZrKWlKwMP/WLI2h6jbY5u6lECA5zsJU8HS+m9ku/vZaK9gaLoyBAg8iyEWGx3kCzPh+l
83MSsfH3eEgzOTsxj1uVISa5vgclK34oE+41L7ey7lQUMbBNIIBBoRn49jhSqGYmihjSsaViJT00
2AgB2DlALfdACn99bKuzCRX4X9LAYFw/Th2t+yofZdcL0Tb5IrfDpNe02wmUe5mUTQKWoOpJEIp4
4Pm3G/LZW2Lp99DmKo9Q53/49aCTx38dG4KUxHkJt8f61uvHDG2xYF3OnqNELQYpx5DD8xlun4O5
yVzLYWf0/NsitCtzQNUSePvzvqR+cjOHz3oMqsRXUJ6fgCz0TonqG7lPpBnD4Pc1ezOxu+DoPVJQ
tbtEMK5cExE0a2X2RG1S8VD5f/7xgqEbzMvdZNtfFAK+bDAGrNbu1OYqhhByapAcc+X9nasGn+vv
fM1AJt63W+hn19GKBmrkLD+FzatXZz6XKLBpM9Idryk0e6LrMAuWs/voLPFLmyikr4ZywUoACq0w
woh7MrLl+0tHMeUoEqbNSMjEJbeBCBZ0lkbUNZ+QnRVMyTA7c6dLkfCYbW7bBCyvbdmC6NiUcpDB
n3+3p4rgjsN9SzIf7ig1hziTI+GcivUNBa3GsrRWGUCJ0devYbeogPmFGAEEkrdzsYnk7JTbOFsw
c5zKAsr4djc2BFWRQquFn9Y6FQQnkcwMc/lIhG+ZtFtNm7VeonUIBXgSZa0E8i5h1Udp2AdA9Nhg
wkdluUZk/XbG88Q2qKN4ErHptWiAzDvi60VB6GRZHvMLCM58k/01agjwEh2XwGK4inldqt4qB/AJ
rZdP73IQQG54EmtE9hCqV6qYoSaxJDmm0ePSlrYec5x9Mn6HZyCwyklJlwWgkPgOoY8A0tdqvJfj
mHOjp4s696I4a4OdBpknhD/YocejaVKdo2uOs8vw0Rh3E230x+0ZcVT2HJ+pjNxnJAjsMXAvKspP
A58ikBXgaZBXBUiUyo3CJn3MJW77bRdgCctlLYHwbL5+1OJm7sqyW+w1unh04f4ZsWWvl7rEQQ0+
Mj7gM43iIMDaF/odsss+Pffb/02tFDVWsRf9Knkt2wHOwo7aO2q4siIUCAm6LwzoDapSG7FtztPr
YxDYiJ8mc0++JYY8p5PGbslCBGQAnljcpWJM1C9A4Klowlnk4h49DeykpmZC6KxqYQayUYVCp5h6
m8yLhtJROFXGMYh/RRZKkHRwS+t2IUu77QQenzNxmqSDUmX5Oh4yEwxGBRt6xtFy5FxQEZo3QPZO
U8he052HUcSJcvFMa7FU/wl0tehoOYkasOpctItBtJjguxZrbnj78yiTIxgySREM9NNT1pnO582n
ANEvzvEqkw4+nXAFVOGSDh+tHJYqzY35K+NEDEO/vQ4ksX5/r4qSGgjj38j3gbdDXttJiwsDckn4
V/2nKPp7BD2JqitPdGjC4d20FpaJzaS51nfczdoM/EGN7xPONAu+lgTpVvegJOp8FX/W7iSnVjcZ
5SsOlTVPzXGtq0qx2qw6mjPicOm2I2glEQsQ5wH5AddmU5r5haKgqtD8uQcVLy7AFrxDqdEP1mWX
Wn4SiKoyiri7Gq0scrvQ2p3fxDjD/8RSrEyuYc1YeSR6KOQLXvczyPacbzAFTHsk1wHiPHlstE23
62v2HlEt5lzTYXLUm3atDrqEffR69Kys23MrZCpaRoUwVd8A4dTeXnBZUoy+Hn4GBaG9bgKjT5lu
lOVvQgq3rMw/6YBRfjPe/f+/7vPsDfZP1KnN5eSObkLzPJPG0m0DkOf7+r2qraKihjds4m6Owq17
6Zxc6WSXmlrqJgFC98PA7NXshtgQxc7lEbpbA2Ise4VIJuggZo5yVM4fZxJnjdSbG6Ugefpv+omg
ZQspPjkXfZYmRV156Wudv/tdz8i6xt979HByw2fYliYvoTVDgY/gcs51/lpVDZ7Yxx0cPYrWMqiG
YzItP0m0sNJqwSSQZ06Vy2HUBi4620swR6t9wUIS7oDH5phrEyklnqoaT1ODWtBIlOtiA1xh+hYV
qelXYGawZPP83prZBgnIWbv6ntL5Rijt1P9Ekr42FQoerDSOJwSdAtiNg7VAoHm4/OK4ETzdEd3r
OERFvWbul4r4u36JhVBipQe0ksprd1c9EPY5PEsVBLY8BWNeNp53p4VgLz3ym9WwxljKxK1pr3ub
dsO+5+G7+X2hDcij86Fbss7/K8HxyDUgkjc14GCFVEJsDpoUqYzCKpPa1f357Bi5lxE+qJCuMn6N
w79QVCHFxo8fsXKgcCA0ogGwdHWjMFOItUon8F0JJpTulFYUVeGM4Wl2gWlh6MU7PRlSqW2hccw3
6HPaM3HEq54NJE05eUkJeH0kTDuUaRJlhrJei5Kcex6WiXCb87YnGqTzwMcsH2xRaATZH+0nOLOt
iq9OQdWxw6bUrVk4dUTlqDD7qYP/QwohGCWPjEw/lB6nuAmQm6ZFxMMdRRVbSE48971yulLLiHb7
FhLSIqoCMNOxoQFGOAaSWOUew932PwpCU/kPsmLMUHFKw1EOggIOgrCxk+OrQylmdv21P/cErCUV
JSsgoYrWvnL8AC7R3339HLFfqdndxn5fIPdqnPqMvRK3K7tKRXLBs5+bCRuaXh9JZUctn/z1V09n
gKo1nD0oM0rCmhayEQTER6glcZA8ENVi2R7Vr0BEpwBBqsgjMOfwAJ4Sf8F2YYCVdOQQuH0zuY40
0rzvsq+PWEBsbnmNi7JWwdo6ZrwyEghEPZmx4DB6Xaq4940PS8Q+sVIndM9sm0AxFqgasNG+11Vm
e8PdR6s3gjbj3haAUNuWlYGBmH/90TG8vw6wvLt054j3w5YMy2ph3xz8hMJDQIvEyMvhyIOZdggw
hY53FQq0EDnOnAEgLreB7+JcxblU+BrwImvjAEhkhaCjEsu0wgejjYhuEbXGiOZy57s6MyYAYUIm
FsWX+W8XsNI+zxI8OSORhTxAmmhRBD/iN9r4ZYSTt41TznwhTOYLkF21pWmCW+8ZdPt6Cj6FZrK4
F0bJsYgYpRJpz1dpvsAmn6Wwasyx1QE0g0YjSYI5NVyBRxTMAY3KBPMELPTewHUFaNJaCM58303e
e6L0cKmCsipy7xflR7qZcgnXelDbwkHSgENuVj7p40IIOa4KUAmXTPnOhFMIZX3PPhjYFAQTDYlb
nMVo6OmSRODc+MsvWwnQIysLrBPxXRMj36r9PEKfylrrUaxK1cVw+Lb87aJuPjzhBOsHD2WgxQdx
ofHnC8ffNrZlyvQJqgOaEZU6MXaWGdQKvLcZ+Y389AgVErgTlzQgHfS5svwnT1eLdGZLqV4neL1Z
5n+iVS494mmQzgee/1IeDWGY9oRZ1EBTz2KJUvB2Ij4CJRaecsLp7HLXaqwpvkS6CtGDOfXfnL6R
DEHyA21sUJRo9d7iW52wRBxas0jvlIplutGqEW8DqVr90bvmCmgE8Ysmurxb+IU+/vvjbYeYTV+F
pAmTRtWKYcwRtAWw1fh/C6QXCs7WO6LXG1Klu4B9hlByx155nGk6M5gDW8sd1RM8dz90TezL9NR+
rkgo9/cgGYHBCD2dsdFu+DSbrTV1HYEVYT/dns0vUuKWxly5jTOAVgV0yPCk1x8r+QUYDpgIhLdj
cvMwMVdbvEDIr2aG1m4BFXYYMgrnKKydG6OZ3C9z8Fi2nytYZ+jEA+Ajkd7PZnseCC1Z/qCHTc19
dr7WMTsRlYtNjDgf8WcOyP+iFZSZ/mnkYgHDRHl/kF/qlI3Kpoyvq5hzh+RiuHTR6jWFMc5TE9l6
0oDEOeIj9kX1JSnv16+22O/LvfxYDB5KwASfCCKkGC/17bgQJatzaGbJTEMt/oGYZBa981UnMc2T
U/oymJAppQVpsL7xwnvlX5wzPoLDZiHTVt9DznX0hIe4UUcnZiTlZzvgzG02sl1MrClYB0Eqnr5N
AvpqkplYh2MGyOAOK/XDDblZKBznZ10h2kjNp8+hEdphaL2Nofq9SZrBbMiBnYmzdYni7mdnkgGF
hdQzis/WuYbt68+gdswIOBUypUMqfcQ6TCFFoI09G5LutAG8HymA35+Q6xzZktzaeDCM9KeYAk1M
Czawhbm206dgn9CBhLdSMO8DL1fgd1HIxfLwS8QvRoWI6HoGMH4qh7UdLIfdSFCxSjiFs1WIFoc2
qKfDIQKgb92WuDxnng8UrUErYEFjdVKeJ6VvWqRZWEGTTt2hTMaHmQK33K31QoQzM9BYuCkrDfXI
eUiut/XTqrsK4qtqud39n0FGmQuS53hJbY/XaWSMGDe5rxIUlwQsVROyNnsJC6NR14UJRd6stAKK
4xyfcVmoEqNhz+TSTHNuU8e3FdctfMjn3v+0FAxQQEn+Iq3r8umT8Jw3T3FfhWGg9tqNpFONqqoV
rS+70+Q+6xDSdPUMRinDmKNP0bDDgN/fL5Ku8g4t/CH6u1twAsvMEHHUQ429c9mW86JhVkSRDbVy
CmKVq4FLmE6yRgAd/wRFO2VZE4j+fejLBdpf+bMHSkYj5aDkj/Innw0uttIAblf8q3eRf7uwrJNw
GHqOXdPvBDZNqdBHGtqrnIoJLp1BOy8NoJuoWWMHvyY5zNnt6jR7bTdB7ejkipnn/hIZvqMcyQmx
e7xi0EjEIOWJAiETHWkmYbUHjKFaZnn7D/xyc8m9XA+DKGFMR4k+2KSF0r846QaVFfkr7l/+n6w3
NFTo37qnaIxgztMGZWC1UDzz3BR+lgmkaWnwAyHzioIa6DU6yKqjFHhBaw1Uf+N9kp1AXMW6h29f
5sFUyjop0IRvgAJeeuUlWCIQs/lJOh7zisaK8DjVD4Q9iTKcpUe+18bBjwoeD6jSWHuYhRhAD1Yt
/ZNfpuEGQUbxnTTjggj/JJNBYNpuTzPMeU2u/py1CMuKFE2wPQ5PBwj7G54p6EZNph47Z2GpdR1S
qFXgfoxNDDGF+BLOSYJ3PhY3a73liN8bfUhVvBOmegrPJn00VNb/7uwUMwvKbtWAW3mjI3/eJWby
mVos6rXhUoJMfirB138UKwxYyiWI35l7Z9AD3zabSY9Ye/PvUGjrqYfrYjYDllyk8CeDwBKXi+60
2JpPrZp0ZavvZ0knM3gOXoxTuk86Fugac7mB80gO6gQiBwCfoiE1A2NK9jeeU3w8aL2NdfvH5kG6
mP61tPIxz2ioZAfW9l9JfvYk/y0hS+OBtyQSRcQsWI5O12NbTVbWfht024ZTYMqncvbJXqyCLSGJ
7oeZPdhEiKPawLsWL/dG3Y5V2L3ay2pZtfoozhN6v9qAHiRQOXZXBtxXiwEYDbTVGwtBt5GB1Rdr
NnBQPUIACKYtnHT+QPqWtxQ8FeooyukxTF2375K2rWSZjVi+fjTwYnQJepavojhKmmK65Fy2knY/
x+xDshC3PNp0E8Qhz0DRYgaOcaMl+esfRg9dCf9x+gHneIl5n85MGpKRmb8zYFVqS6R9n63NinmY
jyyx+cV3X1n8CZfE6C5onT/ejV0fddGl8lo9zVbO/fvmqdm9KbaqMwoCggNKX0Q+IxwTKmM6F2IO
yzw5LqIGEc3DB1PuKiiyyv5Z/L+T/w8MRDa1XdhM3hJU28t2l5x5YVL06AJm8bFtYOIIbm06Z4JY
mAMAIL7xc3mzJMClMfd9geZY61/gcXxDLd8AKki43IdV638lZDzW+1wczmNdAgqjK1J2Md7BstA8
7VcPaql6KqF19KwyAih3U1eTwQA57064jxFaMJ2H3qDMPcgSP1E9FY05r+wbFvIQSqBqrZB5rDwG
RjW85zNwrILJDfX50IXHphhIaLVtnKlxZ100PfI6aAUll56ccWqrrUAPIiFpGnaOcI3N+I/ioZ1v
NSziY29n5KOvUze0rNZfmga7R46VVSAeoP9nf8XPigduvDLsc+jHFNc/QWsKePWXASjhNtJXUOkr
BhfyccDpUtx74arQ57o/IeAO85nR9jFWNCiVaSgfJfqySbweFwswOVGeCgX587zc64pb7dZ/4IiD
46VpttfmZsXiU3jc5ITkW106jRq/+GJWLU9ac4G8qq4NHxxspVg5gBI+8DWAc830m5pihO31VAZr
zecTw1FJMkflxDGRJ9f7imsCCw5Q2p0gb/JxurzkvtTUfU4M5e1rXMFa7Y2SQ8I/i3/+6y/TLX6Q
T4GX6fn8lHkMCyYRkCT5AsPzn+FOk7M4hfMGnt1Fx5otfneBGTDA+4NcDAvQPieVfBoAIrqyFbWe
Si8YRieONi/RPX2yEPsOko65Uien/thQL7/RVF+bOwMc67c7Kl/aTK5PDw15m36mLyvKdTiHpJDJ
kpohFY9lmXTjPzX7wvyeSVr1dLqjd5mr4WhP2mQnXcWTaz/CQh26eLrbC/8BHxpsIjT7ng6Aa1Nn
JmBPdqyjvZhc8+hDhV1SZDBacoZ/ZVYcGUUkP0EjmYE+a6miK56ALmXvvDEkuTMRDx+2HrWvFX3s
PkjAsOuvV6h9cwhgidUFOWE7risKSkXFBz/3GYIK6BpvOmoOQfKX0Fdkz26d8P/Ldl3/1/MFOFSA
SaFhP33HUNgufCcfvWOWFmm9itKCeE14yIIVOzlzeLz8CVGo59DggTf9XOOGIG9e0cWNUnJy8yks
OW1h0IUGAeNmy2HdmgKO6Nxc9PRw3Owmg91WMxsZ4P+0A2ukRULiOoGooMwdVnHmDPzSTuZB+a7O
7lK0GX3u6UeitN4s834xNmmreSDU0mLPcNLf0KsL+GFzwrJTjo6sXmnwTqTCYHxIfCIRwGSwQyWw
SirnmAukV5Fc6U+09NKm201gnnpMtaQJji6rpheFmNJXPdsGw/OXEZKjkAXW494GkKZ3rYGrBwJz
5CrTulEzt4DKnqD8iGTPoDWK4p0KrvIXq+I3+UsExBagUXVDxQOhnuEcmYJ/+FU5i3yssFjIwJNH
F17A2iJu+LX8ev4VgF43N+glWJ0lhi3SrZsPzcU0xpH6i1di/a0pIC4irCGiYHSvmGw/wJs95I1Q
BA2bSBPP3FOSrJpktZ/kniK4jVQ2WM6gKsnlpEaiHw5gEvP6szcJnyiRyJSBFMFdYkZdsZ6/7o+P
gN2nTKSzocZ8g0KGUKREtEcwtlUsC8KBjFJ7HAowB+EnunETSIjO/P7LTJynSqpbs7z+zRKbgnbX
pRKEikiEV2gf/mrFTYnnc71tBctf6A4CGt94WQ+Kx5r+crhc0wbnPSGsjAFIDlE8SIKJkHNfEzug
1r6BJBwPSTF9Z2EUMSZgKJfzNtF9SjQKrFULh67RDnfTeGCgxFLhrqG1FimIOAsJdAAeU+MLfNCi
ynJfCcpSvi/cQSE68Z+E24sxeE87zzOdBAENC85EredS07qL/X6w8EsQrAfq5AqkkVmgIp64i9Kc
HWpf7qKjpSGO3qaI4kEtfMYJDEJhUg/H2XEue43o7ey99f9F40hjvv4jcx7b2cuaBJzAQ3dm0PvU
x9UfL8de7pVYStUZNR2J04RKny/UtXUUTX6J/UPWOHKyMFnY/BNwHuCNJV4ZCy1aFDxo/Yex1phF
PyqHUU7WxhihBtaAYDbUXdwFlWjopqOA3pk1mWb2k/m8bByNuNbCplmw0ZIRjvivrYcaNsKS/Poe
qNFDdh8gTqz8+HKAV83zuONenR3IGE/1mxPSb63QzPsgMM5+oZ3Kok/r/mPILzSTHecmIwfl0vhl
e3/qtvOWLzyqIYryjQN8KtU85B+uhVM1dIMrs1kW4y+bEeR8VJlXl8fOZqXkEzvML26X3tn9+VUo
KGrDLpyOVI6TZasWBNz7JuTRIuuqKlXaSLWixR7tOnawKzrEXVD1+bmT1stzJQKjIIbchDinEndS
kyB+/n3A9oFkM4ejr5ntU/WfDjZ8aQRwR/RlQ0XrL6fCkxY37bZ1+euhn9hQfbibL7KS/NLx1xyc
u4JuOT3L9fSpsqVljB6ipXzX0H3hbyeHPUOlNeml+2klZrWUt0XbpS2gMru2PaRWYNC1FICpOAR6
gy9MRrVTv2CenrAUIHs1oGQ9krnhZvnwHAytNVEgQjHfiZIbYmU4QMScqtVhU0Qg7S5whYsy62ZX
RtTGCMqgiotDbNyFr8zYGESTeoRQz4+1R6m60GEUuXI3fgyYsAQk9At4t4F1Gp/5FWJX/NrAn4tB
+VWuHGj5xihoCo/pGPO9K+tm5VV4YrQLzVklDryZtS2UOUnHGq0865xn2R8WQhWgTdOqN6dI47hg
5SWSlL3pxBAVy+nxz6mNwapwPu6qi2rlpOZ5ew4ALv4/87D5Aex373WpbrQNV44aOkS0D2ZniEsZ
8gxMZGI9uJWtb5qudfiMEsmJm7j8oX7Z+kZ4ACH0a79PE2KJfMSVSQyu1NjUje2TYf2ISEBxk/P7
ZL4kYRScKFGhqX0C5+R4d9ID19b8MGneEaPOVCJik1f3zM3GHgYwjLR1xix2NGr9ySlFGy9vI8ay
uXMKyK8rN16b1R4BpV4V4hwf81nukeWgLTb6fBRrThOgg4FmKqvHBfrdBFCDnC/aFqAszhTeSwAv
L9GmJI9IYUcaCRcOfcQo1pwaJtx0QKX0QDVMcZhixwOfInpGMZWwpG9fjWW+RhDd+66W9E7VwcLE
7oJiQaOUZ5QCN0J0Gke7M78m4CX8BoVAMTkAxJCaN2kZnJf1OAS5luVI+Ys7LEphkuFGsV00Q/ez
OLmPfZWMXSDDDo/C0hsUBL/hoV2AOkxNzY+ILrDYxoQu3+rs30RpQlR+1k+DR21d7PVsHSL8ObpU
wY/02U7slB79Gqk9h9fv+JAIvFg0ukFA3ej1E4GNbJbD+S/MQmr+8HFDdN/4ej0GdYp3WIV/oT/M
Q763N/cqZ3+Yrf89yJCgTh1NgLF3aru5IhkFl860LrkDFfi1H+66eHrhCUhLUjc1ID7rz7ucvc7o
cjs4a/8kCtbTOnkMp2gKfwKd+nCfvCEcWFLsSAqxQ77na1HTy2nG5AudkBOBWGpNL6U1dTXJlT5t
EhgvPZsh2qVN/rAp7BBBlmXV4KoWuKstaBLMvl4M8fDVukhx4grR87o1thKkZunvHmj9j3YLa+uG
Lm4J+xpFV1WnbfF0nxl1Jtit+ttA7CB6Kb24vPWrh5TJkqgAzMvkS6kqpLRITJ4L6XEsJ+yBKdj3
yMeyr6bReivI7zg9GoAW2TuAG/GssXW6QHWKZ9RhEMmi8lq3rGEfWRXPMb8xJwTg0UQv3SM+tVAp
qGhk9lbCOMVBhSpYnjiN5kYVLmI8nt0ly10KLGa1wrtsDUV4BU+dNk76TF339vz4NpIIsg4C8q6u
beup9vU8hEIXi+80ycEDLYRxGuii/3Gjq3YbLbmt9xf+EhG6gYsrrPXe9VuHV6IXy93lQCtyfHZ0
75ODL98ZaDwnlgzsI8qjm8u2uMj2Ug8/y8DFEqc3c7RHeqVpB/Jpxx7RmXDMaVM74rQGy9bAGR/U
jD5yryjy7dOeTSQ4fx+YZQ3CSZwHGGweFg7Idx80kcYno/+7Spj57u8rvhx39uKMXMgK/Gk0ROaE
QOUuVAjbWuBUV73KHTDlXQHrrSykjlXGUlNJeksw6pfwQg/FQDdPmYMHbRL5zaUc8E1ftDEeJ64L
zE7eqki2sHW8fMV4n79BUjmvIY+q4PfsYhHx2LJs8C/1/3EztmEARHZAoMR3zGyKWv28vVedxCGr
g39mO3rjuk6MYTjvF9DXhhlsGDg8hlP+Nwc2AKZMMrn+/OYRW9rxHHWClmXOVTrV6OAfKJzVUIOz
k/T36L88wKkVjNojRQZ1l+Nmzoouc+ZrnB8UKv0+QSatsup5VpmnMrp1iu6sfjX1pbS6gAiQwyN+
YCPHHBl8Lh3aAwale4rOqhSbBDiDBEnL7nz/k3FbB/VJoMsN591Ockw1jUzXtfbl4qATG87bBbT6
k/+VvmCTdHJOeEgAXPKjjpchW4PlE80zjDVyQolIRvZw+mrb7elB5OKbNcXF+SwB2YTHFCw3VWm4
ShZIiWHgAsZ6lZ5SLjBpIzOSqLFGsEEobDOOirJ6qPrx2tq1cB3vStAVylxIqxel8TOJZ30rj4sc
wfkEpRrNd95B7t3bssjf2mljd9SX0wD3tykQKQ/hcoYmVkjmZlZTaQAAQAx9GJTxYCF0eUbwRkDZ
7AIubzPuvhDeguXZuVFJSXp/g4M+jjsNgqQDQ0vpkFZlRJEMT1WktuBtD66N+Lq6ck3g/tMnLBUd
vYsCvezcsELVQMzwQDNeLUBI1eygKT5dKMjL8ZHt/w1Zj/bY+2osKMBFbxMoQ2ZD5mC1H94HWFMW
Fu3dXoCs6fQRgz77JxQxWrT9bQG9Hx7ccc4Al6PnAlaxUg8duNdKusPJyosGw3UfdmVOWBg+/nVb
mFlmh/hWaO+CTy8YGrFG8c4bYgUABP/VokvxEijhIbOb9KJRK1lrGZVJvdHl9pgDUnSVav9EUmLd
cqXIb94vP4pJzHZD/DVMSo76izynMFy63PoduMBPfdmPg1NZK+0C/Hlv290COdDecnoyQ+W6k+Nn
ZtYOrOI6kX9tE6WbzstrTTPUqCQj3Qsq03I9iQkO20rIXWGY5Gy/aIsa8mMeGPitZ4pV1y1Ue0IW
laCJGbNRZKqLoLmWXlxaocNywhJNY+HX19gA5s3+e97wIzrd6YKxorly6wimXwcvi9noKvV2Pui3
XmAybs8PpvHisx3XzvYny2iJavS4h67QusnuWntlvNH7XKifHNZ6NfUavw2YdKar1JHBF+P5iaq9
J0leidOrtv6j17lqiq3J8Wnnwp1xzAV2u75vof05pJZYspCCA4n0OWuq08dLV2A6NbTd6HFIJbAQ
s3sOcS8bL5AwGp+EReCYskoQtdv3k89W2Hs9M4CJxzmW10x9E0grRWgNye5hCTlxrnpoNe94Wcfa
/WWbrbe1XZxVJuU3fXuUqQCHnGl7jKMLt9pEGJtUxUBo8/4nD/uHCnPlNylayYVP6bMgNgd1+wMm
2/uReBiECVSVI4vWOXw7CdxawQdh/kfFDAfFSCO1Zm5LdLQn57VhegS/9Z2E6uW0AxZqQFmf9TDk
ox3XRraWcy4t4FkmVrYISr2vfF/TDCy39UWz/ifhdKwNE5334U9xVmlvMOJlUoBRGy705RT7NOpH
tBSPxZA57wfCISy/Aqr+aMWtOQI+jUKVDkKPI3tIuGeR6Bv4kvz6prbYYhNizZNBUegrwIyYFQeM
P7J+quY0bS8Nw5foqHFNGhU94FMMwi95+EIbVlv0xJBElb1YlO0DU7XERNdUrocUKjspB+99Kwqk
hRz062eYKiy4+j6/PUwpyCsHrF9p6fqvnSWBzZBfrsubi9oiAu5Zxb+rTxuomCysErseXcUXHtQn
dK8Woha7nNDZ3NdpmXvlUHYjyLSoiL6ogNLgEdiZeX7PwixVi7BFb70/DTYgKuJP2uQKMA6CXUCs
EmeSbN2zpoI2fTe0ipRMS9NNvI7TzOLss5IlRcrO//vBr8BWSro6gyfbCsEnm7spzKPhELBl07iX
x+m5U7GMgUGtk5lcT7tgPzFtQT7JWND+NRVmihZ5glewLB9gMDBZhI+AiFojBEBbdGFK/nS6MB+s
JogSILzW0vx3G2NQxWOM3OEnmHy7E5d/F2WtiCSlJHMdkR4oxUckMAGG5/zeAYPD3Va3S9IgT+Pi
Nda+Z41jrGMaOc42WMWJd7Nwmu6RARy/Ae/Px5KQjkrCO+D2ZO/2rdgj5kN/27+lCEmJBlR5haK1
nf8iLLC5ftEgLo6MTajrdFxTnlNNUVulA6lRC5fBmh0vThWk8GepEhEAgQZrmSa13K8TAgByOL37
43YnYbzdjr8GxbO+aLtC6DHvjTcFEfae0cgRI8KVpUbrlUEa4bkrYpZpwuHGdyrx7z/NIU6fUlzB
kkpEZ3AnM/3wrcZtMJqEl+rxophGDmpCPpKav5kxz66RUeW/eXF+lfufasJNXG0BFt90yG/c0IFe
FdzFCuHPaAW48TFHAn/dJRyzCBdr819OqrbBE70rAOrr4zi9cvDWe5TaL9JmONE0Odoq6Nhj31Ze
pNyU+O+fgz2zjLd+73CMqASdO9QgMzlp6TyoVour5pfcA+Qt1IHUGcgJ7/gGqUk/FUO6vilhlse4
DFDG5yep83wJ4rBbmSCa9ZfwAxk1hCkc4fsKQEgl8MBlohgKNK7AoGuA0nOJ32j93N9iXz6DIYS8
fbdGWW9XH6CuDsOH5J3Bz7N78NcVBzqaT9DRygGXaw0HGESK3F1K52m/3LAlhln8tRI9Cb+UVyZZ
+Saginms0yM2wNExDDlfwyXk0DwP+JqSvbgh4ub/lki1q6ID9xArsI0P144eJDvmeH8SNehjUYLa
iHbvk1lN79kaBvvXRIfNpTmglUOUhmLZyXBl357G9rJOoXEbzxWDoiuESiPOZlpeqaonNtn8u5vN
IjSCz5aaj9UdDEznTLHSkJY8+gk/W1AZDB1ngEA4onQ8Cc3YSGo+6tA0X6WMk2TjbLex3pX7ROdt
Tj8ce1P5syM8SaVQhiKn7WKD7RfLEoS2mJf6W6BQIles7BBtT6CNsnlagl+iXkE9zdEg81OV02N5
71b4rZiqaPZieUIcmSRVRy/wRUtrSfUagqlQvsrVPukWaXJt4NSK6BNNfbBOm+o1NK7IWtfX0s0o
/lcD1cgC6l7AWVTb/du5fDY3Uz32uyElCKfrdX2g8EqTOyLIzZ8+Tizk9zVh0Ikd+OYy6bbWoRFA
3jpQRy7QGHeVgqG0n1Mh0sO57f0CzzmxgnEsoB3DFP01GYs/4jDTAz+O8nXxzK3PI7qKqPVrIlKU
68lmP4r3cTsMurWW1X0TOCMCjrWQ84q2bhbXIgC+KiWeB2wCydxLUu5yPjHEnVja0pNAPCsOtPCv
WDWoY3crR/IubCd45RmbkiwNb1OuFNG3rHz3M48y/8w/LuW00k30me8kSguGFt28dpK8A6dOb+j8
5Xyf4uV3aFlsXLPC59WOZNkpRh2rwAclJjSUgjkZCx3iEYr0V9fA4dEJF4Z/jv0FWAoMRFAuaw9w
IzkkXw9+PLZ7GTMIg+3ocmhk9+HGOXRi4xJuudcaOuq1Bd5fdwNoWjk9SFirqji2NuUm6jTlRh/s
cNG7+rjmNbECLxCjYmHD9GzfvC/alncOWwDdCcMTKAfCt/aICEduzTEgsiDKYG/NXWk1cdBLDYcf
5NO853YOKxBKocAvsVfmowmF3fPkbkofb9hgFnByHZo2TMoWdgXk5l+6y20eMQFMloTyRBiT7cif
izxl0K4y+t22YXpU/YdnFKpwenoRJ3xTWVG64OIz4sTMVE5zLp3B6fK8FktQ5fQVjGRxTfKNMf14
0epW6MIkonS97WecwmWcYirsxrT3uXEriu8RuyY63AJUrtbCs2JDFSzwgF+gqP+mWcnt4Zyxtjqu
/MOWaQ4RbublN/gblPPWWS5ML9uYyyWKZF1JGMltqu8hBcWXQgv7B2aQQ4F2iWPlIiumTPzp6tdW
Kq+I1QsdJcS/8NJJKivBygTg/bJb3APG8pO9MxhvX+qnN3is1e30GiYeSh3dWUe+sFg7DpIQ/rIy
j8m2IngX35fdtiEZqkk4sgrU+6qPb5bW3olLkzGt0uqpQAHm39/dFKNgGQW0wvLH5ygwspRFQb12
KeovEZhqYKnY29/iQgGN19qEZzHd4W1G7OmGF/hDcag0uRrDhU3eupIylT1/ZGWaSekXMz3i5Sjq
aS1UVjLy4Gm5z0IkIO76JKYpf8ItjfExdStQun+8413yBRAhsq/X4E9qblGWEKi8FBwBy9yjqUa4
lHrYgMI7auhT3zVsBVzsiqVMgyxmYn+uq+6kw22bdoZY71FGBWKxOXHrYdFU6VUAtl+ofswe8WXY
zdLj4humrufFI7PxEG/pWiBpOJOYwvRjiF6TWtwIRtavNHDJ0agqSMyH4ppX03hp41HAhWidcMaO
G7XqQ2G6VX3pOkbMek0cLKYIDCkKAmmNVH0C51tMm9Kx2FlPkr+1xPhGTwlFWVySjKYr1zlbeAlh
wePU+jNapMNKnQcO/bFNIGFItD13NstslTNaDRlX7Daa4vZq/OcZngNdprYmEFxs0k2cVDSWeUWQ
ViU4qF54BeteTjgedMQ7/P9HBGiopGUJl2LWDgz/sgQANh0umU6Ky1/Fla5wDjK45JirgxC5mSXC
CP00aQ8OkJHTzW89fob7/lCoo4NmamRIWtUQNVHnYq5+U+94q++YGMoRPCmPm2uzn7lBVIqrDy34
3IUWq9UgQkiInX3tpUFhXVo1pm+IcmWfcyXDwpNtP+AtNIrlM+dq0tRT4zDjPFfv626HCDjYNKO6
lgpR4ZA7uztEe8e8RH766MXj6GABE5IuFwXYRvDfxPveb/9c1CzTIsXQjMS13qlaHdMWqYdn7hn4
4Q675PSFpWHOBodDHB/SpKDLiCkhh9SViIx6AjTcygiFNCLbAuLFKaXLuWjddJGeB7Cn3gDAAgeA
XkxMtOuICx8TDuVxlLJFgTbAuDWxM9RkJQ8iDBQycR9wWVyy5CBxt3/eKE+RjRt4043QLOD08oYH
I3LMOU56CeQWGNcCGeyfvCezCO/n5GK5Iz7OfzbG+Yrxpjs4BkxsLaXRHs3x+atf9VqH3BdtSC/k
zDD1RqAEMMmvOkHIeVMcIvSSAWB1Jd70dk5FsAkVqZjJS6K7VXLGK1sqW4CdePgkVMTokNZEhDFo
1CiEu6zuRvB9RIG11gwwFU4PDziiQzzwXrns7WWBY24INJfKISUqiReTia8MKsRVQcKi8hRPnWdH
53tzVE4FFQJxepYxXkHGr2oonYD5GWDyKxPqLn8YsY7Il0L/MQxykcbTWFw7zkZeTZcvM6ZnVfLZ
IHvIJskIc0QmvDdBE6D9qWEdD3fKpfMPXnx6HB1xrVdr7upPUYkf/QVWUbPmTVLGPhyNg5FH/nz4
TRLxP0PKmlsoszWKe90Zh2dpvfM0PgNootcHuIDogQgo7hO+AYmy2u242whPWpbGtYFWJ5neQLzO
VrUJfSRSt8WUEVjYKYBY8RxDqLtvFqOAy7hC9MnrvqaYyLr/Wt6djVa8Yg8gQR/L44jD3S7qwH8+
NGOQETgncmHY7fjdC2/X90NQAK4ujhnRyR2DxZTWH87ZlG1aex3lS7IJ79l9prnvB1E6XO3HkKJh
Z8KHQoVHkVkYDL8huc6EJKRVoY1j+t3kXfpzi0IOaWPCu+N8YL2tV5HeK3zYb0TXUF7Z3Y27yN9e
GfFp7/N2f4EfTEujKugr1dSYf281rVi1xqworIibvwNuNdxDZUo7e4lSAOAou/1dZNru5ye14f9O
HH9Ikll0UGPxiUBYwjXXsZm9ZjdVCQjG3pZrO3LBWX/I7Y5geHf+Cbp7pnXfDNzeG4ppRi3jyg4o
XeWOWu4f/sdTiPmQhb5pp22bQQl4r3HmboplQ3EQanCKmQThvY/rpS63yoi5Z4fAD1AqTTndaei4
AkcBayUwcM/SQMjM3H0Yi6glBtAv3JNEDXwlrkFtKapeJWUcV2xYYAKVqmSeLSr/6k1Q+ymIHgVw
lmJREafDUfHQFvPxOb3skQP7OTOrll3z1o99qxhP4FopuFXgpeqRwOvcvVSqkWOsDQDfJI+ZLFdF
+dwFrDsycHVML/lXriDJhYGSEhrPrBCjifpgyavNs+qoFSMG8USSfxE9WRNBFAUYtrKu5md8gq95
W+KRpm7e7oDoV22NJM3VNgvcwYqXOBQBCD7N1DTsoiCYA1CXGIkB6V3GS5KhEDTDMbP0UTBoWvaq
NbgCkGpSLBoPKOJR8F1ZDsQgQOCDzhKfVq93vJuFyYY5T6u/aav4t4PjB7gIjJRHT0Le620Y+Zm/
O/Z9jYhkquXcopLT36/7q/yChELcU+nNlVRQ/7OtohZKVd0LKDKF3OLVpc2khNgY53z7ful/Jcsy
2iyFUmIwlY2wPuh6wGG/9TCf79+ihzhO/U6fRrp2Dwq+S3NGokf6hsUWsrMOGdPCo1kh4XbLaUr+
q/YhoXDnDo73Kf20bdGuqWXmTMS64oUSpCkuAva1xlmSaS6fQjoXRdYoeh9HcQS2tablI+fAaDyj
GuNMz0D1mx3mC0rfm800BL6thsNtaUIutgCKOYWHAQcAAGuhFPobbWD6y8cpCOgdGSMO6MDAh4mO
DYffMpIL49Swi5pDNrY+OUEsg5XNvO4+iEAx4oUpR5ErRgShxsVqqI/5YYyq2F4ScQCqqeiizUss
STO4K7qZ51a+KeWu5YquAbASF0SxauwT9XQpe36N6HNGVBLtfSmHQEMGsIdncLHbsbynGbhyPvPt
UxLNl+MNP//EDUt5o8DE+ab18bI1D1TjBCRRU/H2cr09tPLsaeVaBgClJfrVI7GXwArPlQU7sO/r
rSdxiCGaoREfJpGBoDkvUQ60SQKbDslpBkTG4G2+gJOGW3OQCrXff+6pBiqGwulHbL74DEpj7hdu
jfzWG1JlmwowGTQf6+fqtefK2XeYEm1AATwdD7dkEZy5n9JbXvcZqI0M/Bslon30tx45JZnsbqQF
OeklM9YpvdSQ7QnUf+q/TRD/a1UhN/ck0AhoIiz3cdUJ1jYcXQNAv10f5NO61x4uaEzx+lH7BRFp
YZvAFs39vkvaEDIkf0554sfiBiD2mwflSZCJNHLaaOxDMwfT2RPV79hAXivDFDUnGofrPB2KA2yo
oNgCPHjo30YlTL6nhcVutXBKdH5PA4/9APobEi9IlrcnwSJi8OWeqo6nKAAwm91YjAVrEpT8gv9H
YIWG1hgkVRlXDf4ztmEQep/Udlg3orH3UW8kuVcz0S7IdF/SANNKDVH9vKHBZ5Cz2EqZie7c0c75
7U5mBV4vjq+9uCEe24LbAElsVMNZf6M6f4y94az47VM14t7VNxt5J+msrRendt0/FSc/BvXGuDMt
D/BtUVYWC0VFYLjJKEYPiR0lCWt/mszhD7ArOFRV6lOqZtrQmVGz4Li03i83NPAWzHrltkEcg5Jn
oHM1ieJagYui8xfWJlvx9WGp0Kt/EWK8KGpLqGzyfvdMSAOKmhMe3V23aIBS41CJwJ77A0BA6/qZ
qG7RsLZJ/NWcMiLaYn7iPQIpsY4vU3odhKExpMLNMBzdDniSV3VvTyYcjwzPIi7mKylbMZPneH+P
jSdtfSp9pobZ/0uTlIvOuszhpS9tPO6RltaFj31qkg0jsQQhqe4BA+zyIt3Qku+KmKp1oyNeLleq
TpYZrj0JCd+DJbQ8BO+4B+p73TLaUJumr7RKzN3bPWhlu5uYuVnvkc9ZZPAjVou1zu3TrSR6jph9
blmBzpTj6yXHfkpRU0ximHbb6O+5wXoFcvzeqiqGf2Pf8qQ7GzLfzZQJ9mxSW8jyHYA51PvF1mZE
xHDar0DR1NAm33yg+3TVRM6icjaffE/Shk3v5ISqEQ39bZlb1soUrIvcv1PAlVZa8PurW4yE0D8r
ADGpqcqBrySXfz6st0QCUwPjDRFP9w5IGm8CKbkX35HrR6dy/lWf/AqWqMAsAKSn041Do0/XIm2s
li+FkGGCFe3xSuctHi8Iq7lh2UV+2xTsy2xBri3yudW+eqjB6tQ1qgR4qSCvg7GbkkDXJZcGJboX
8GPquq3t/Nq5vo7dO/5/HPcfb6FQJpu+Iv5LcY6u39KNhJtJeNugGQqBgBZQMjhUsM5nl4rTvCxU
OdQmgXfrUngYMETwVnmQhAIeiN5Vcn9wf5dmR+nieaIfUKgAb/rzXnfug3Z6Ss+GT6GyqqMa6EJ2
oDsZ4K8o2BvIET3y/5+SrW8ndoBh2tsnIfalS1owXsy7GC0NPsR0Oq1MlwF3ymaSb1WZYrl409F9
atM0QJ/owQhiiMvjvia1msH9yMdh1KeZY9eWOHp9ImTroBDJrshn50d+5m+x260m6ub2yo7Q+kSH
CFMxXmy3PwvZURGQqhHPpGadebZDbsEJ7W6xeKT86fK5ryhVTYUWBN3o0ybnfAtmMFeKBhhA2mki
xkYdNWTeFipHKg0E8rfz/HsYbLemjDd2tVMYrgdMm5rG0mr3e0NyAQutAcET16gzYGdPxTfZAO8H
SO6qbgwKftxnXJazcJ7zbOI2S0A4qWfFoRh4enjo5Fh1wqmQPjfE/+OrO/5wbX2XJWf6KrKpVOvj
nzqudKziboi4nW3DpaTMyX4v3rWDhFm8bWAU401y4ntF5IcNQHHHfCYGlfXj5DDxKjOONvhJhzBR
lCCadKaarPp4uENC9iQI/WxWnu5mWoa2Ez58VjydzPJq7+/kcrqGNcBcKiPGCcfOUm5IR2D5gX2s
3Q3m8qw33nD41R9wEu2zu+ZY6zo/Q3DoZJIPO24ohq3yocBlISTs3LHZVshow814GOE60vgo95+N
M2UcCUP3X3JMSHXlGE1mEDD+G4KtiwfMdelQJ/kjoKmsltknS74Zacp9/nJI9cBl1hvdg2KbxXLH
JhDLztGjUNqNzrJZYLKTp3yCJxsuTrTkQPPXHHXh+RadOkq07QStMFXQYlDt307hqQmzKJ6z7g0Y
k/ilyc1d0tGMs4bK0u5mSMOTDOtLBPKb4MnMSMesJ2FgCAoxUFprwrC1gBdLsRH0eBBN2Uj+0E3J
BFb20Mfbh450bJ0b3Sonr011tdJAEorzAH3gZ1j7nN+6dazrou7rfkIYpLW/RAe2c2mEyVsugkcK
6iOsxkKcGF4Qu6JGOSq31bNo9hY30ECZheqwUq0uNHb3QtatwqPWP0rqR0Q68HadcCsayGSdL43M
V5hfQS+j7ud1Fp/7h6GYx7G/gw4alHV2uXce1Cw5SMB54ifPk0sHjdsxAT6xq62zcjxaLKBIJKb4
oS4yHtRq3Hd0gl4hzbuioUlVUDHKa0zbm/3Z1jQZwWEaSrdtMDCqxbKTNuUOyaLzteNzXwMCvxHT
CLUCy8FDAIRNEGbxy/pZc3aJFrnKU+QToWlnDcxxq6fOJKrclPbKXztvzl0zG3+GBgF/Y5r0f16g
iykc366KMRirbwa1nHgab1YhjSukTDjrIvlHRXMRn/nLz8TNkRSIr09XuLlQCyTFzyB5sEjc5Km7
ZoINv6TmlcFALbmjcw2w0dIbK3AtCF3FwP0CxN+0Ad7dwKXrIcoUZxYR1MwC+BuK/t774ZY3cXT3
I0ENAew0rqWehvVDz6b0GJi9XgL/t8JhfLS9+WuOaiL4KX0ziIP3FuIr0BIcUU3qTG6F51zPBkl6
hMdCpF/NLPvi6JtfcMafMFYwrIu3HsSgzYjZeshVuizB5XhLj1NBhCuyaLvsyFpQDOhkK5bV9DIA
vgJEPU67nvwF17p4EamvfyFQfjIZytrBfuVj0vNBmQNIjSiZn3ZlG3aHHKG+JUU5QI6zz737aEmk
rcAadbNmNkL6WdqY2Y9zyuOnjAupWa0x+AdGctS9DXKZTR1fzZe6S1jIzYeFRR4K5dRBRVlbXBwt
EhBD050zbHA3rVRM6N/fvvBG508F7N5IOBmtHnYLe7A9hr0ML+G3Hw+nqQSCW/dhRa1bpKl4XDNY
+HX4EFNx40gkwdA/iMTv+YHPhzNkj1ciV4a0xN6mwB1wwSJ9c4FT5AHswy9swHLn8vro3lASJsQa
AVruDxEe2I0Nb0Kw7Lyoqhk8o9kdCejvqxAPVSfbu+xXvPFbybwPUICBa8PzX/wrSM1FW1VZLMgJ
8co6ie0INTcJerXywX/JZXpqABW0hcJgtOpcPJB9KF3VaHIncURCs/fxFXZVpevDscj3fp0vzFPG
i/bMnfI+LjA4altiIT9sLjigZ8wgUQW14iEN2a/h+9IpLxzf+RW9YUATj3SWZvqF1kbE8iL9ueIY
ikxNAy0mKT8q/aOY5IQG5LWMiEddH/WOMZz2Tb/Xsrlzv5d3gGzSI3QbnJP1alGZsYCTM7ZK+cr5
V/HrQ1clP2p/nlvfU2/Ca59+j61NwWPA0tS0aOz4HKMDIPggdC2fO8wS308DcdHzLq1GZH0DUAYB
k28bHhRjqubKOj1MmJlmSfWHZNyIuknHCtcE7rx1c3R0x2aLsceMzlAyPnNih9++PR+GZvBdeQGF
oMLB/MjR5Jf05/N+rA6m0NUCrEaqNJDLsZhtjskW+xDaE1YMi36/Oi4v5P+E2yAQVSb0m+NhStAq
FKN8tTeYXV7flREhvwlecp7MG2YTMF7GwbHE8U8gcpCjuRrb/qpMMOg7OPg8f0qOLkZiqsTQlVxa
97AD0E70Wspy2kUiI6GtXqbw6YNGtyy+TGPtmQ3rwjXLKksoZi9oTNws2UvWHg8aoQP99Rmsfg0D
Z/RtGFVLAXEzeYjBWYnSzfkA0S83yeipZgpd+/P48iYvdxCJ9baAvbnF7GW2G5ydcPiztG1gxm6R
kNaO78TDaFfezEHmNrjJWJygQuWL75yabeFMABmhmeSHujSX8b5YuA+548PiFkmkdNmU3X0sci5p
dZs6Xvk9khXhLRoiOqS9UbNS8rEOT00yZitbzDMsOmtgvZxKUClVRTQum0gWcyN8L0xOAelYXylV
Yhlss2vmk3N5Fxi/XO3xj6wSbQuIMH7U0cJaeOVgvZ8hanvm4E8nIb7Vgt/WqmxUfUr4YB+RZTat
C7OEq5dsEvmWH+AKU1k7m7fAAROcu73BIZy+NYm1v+2nu+Zg1HXJi6a0l27HTGx8LmlfoVOfA0My
iyGQgvxLOABIGE2pM2GdU5GyKzNNbKhDxdCXnf1Qz2AHrABr6dhwFcNgjYtfDAa5HF7GoUBi27tg
6UUb0VGNQFZclj8yPcYcH5Nq1NLZucQZhKoDW52zqSV3z8oSEOU3zIpWHb70wh0nQJBXGBV26HKi
H2RMLwXvBVA1CS3cNlZvwEYwwtzIUOe0EGWvqJWQ1sStcAe5gjfxlLiN9rnOdR1LvfkMvJZgll48
SKpRsg1yP/WvQZeuBReAzyKJ8C4hI0bXIPXRr62JZsWbYoAIHcahAJlbcPLnv4LuqW/RgWA02f4J
zZHRn0p0qA8G7/OS0XcfPq6aXuhWNZkmBaWaJGHx2sajOJhFsshdriWNuY90M1+tYGmiJctlLe9F
qZYMmr2yTg1YGW3pS/Kbg1TR7O5AyQfxnBTSjF/6XVHDvzYFtxBYg3vlLtqhxCFBqSvB7Pnr/V9t
Lg8/X3ZbCsVQ/7cXPgr/Q6t1SR7oz5baEVAF622eBPu+OB4rvJ4bbipB7zW3mdL2ReZGvBCfwKjP
TJ+Nfz+zrKmiK5U9Audykz4ZlygKdkr1YYu5lKx7hRilTiZSwT0FkCXSbiULUrUDphRx5S3zAAJC
k5xHUIM9SWhvK45Oqfjp4tjJxNP5Cto6rblkXYZW8vhigLHIKCyh05tpwCucQNiAeDp3JZyS1bH8
tJICa7l5diF7uk7tJlygpsOiRzdD7BY3qOROyBigwSMBze4AELyHQMoobpqylbsFKr9LxlBz3dc8
34yjrkPFxkB+VhxYm0j/DIYID95cMbRSyodwKQtpEeho7+GWu/tLPjkmqz3SvwzqVPhU7ZizCeeg
9napnuV9wX5CD/iUOcNNfGjJcIA77eGzU+iTDLZcKO9T3l7oxQtBXyv2lY7IkN286Hw5d8WViJ1G
zfrfrns3JGj/wihvEdyDMFo5QHS4Q/jpsA+r6HTEAGb+6cQKkScmj5FlWVYiOvU3jPJVuqLiQ5J4
SQPE53pwC/Pix2FZOwUal7oz9lbfWng1kbYB8wSZSJipkL+f06NARDsiX2ezsY+iAWZrsmHVWbgc
bsfcLEQIk9tljipNBd4REOCTVrJYLnrEhVX8BUX6YBHvo1mN4wXCH5cRio6Y+fLogoRWwLsKv21p
5pmxhqlBlRRO2hNC9USHPcsH/xaqN0o9VWfMzQGu+3VH+YwdaFsD/BmIXhxQ1HEqXnx/eZ2RTr1g
SQdmHKhLBLYyR952QdPAAkoB4NnMtk//ccRiMIc61Z+ChSdMe6G0PQWsyJx6pFkEU2Hy4DmePTX0
1cUBfGqQvmWg+l1GFH+ef1PqDD8kIqCggqjiu6cAcZ9pe4xTJnt6BDLKLfnzqvsbwPJmH29u0qvg
8ueIQNUGRfcuGxjQ6AezmSQIFa8CQcrwd4ziYvFiWj6WSPqo8I4JRW67vfNw4QwbKIH7VbicbaaH
X26Jz5fUDjWos3n/Gd2qkkwlanltM+CO+p6IpQtB5L4lrs1h/KIvdPftt/Sh22/0/0YakzzggEA/
l5KN7unRrnupccUol4Tq/OravINlLY2K6a+k0rTiVpu5bIG7x0o1wEeQ3mkzFb4GX53MJiyDXyfq
0/HGgxu4VaqyJyOdTp6gXy9uhZE5DgSy49P3kkg1g8a2sdVxs0dacWqYR90h0vUng6+p0ypLF4A6
xnrsoJVh101/f9O5bv77wQHOAu2zpK4GSMrGLIy15c7Swn9KxKEt/8OvyIrfMlxBooI26tB8aX0m
Hjl39DqvRxM3kANKSD72P7SkukvtoErkUZNhPqe4bar3CIIf0QpTh/KjXQpsH8F2yGU56dy86tCT
9bet2ailRJA6jiDqppSUK0Spi1doq7tBXvmZQYlmk4tjEdDVB7PNhXKLL+kv++nWY2zmhx7SsZZL
61STEcGVHx0YXxMi8j+vmHuT5fERRnPqPY0ZGJobo/ZdMLeMJgmQnUOzMDApNc0fNDl7Fb7TwCEd
shtW/E4qHxKb/U6XlXrTKOzNMPQCStHZ9ZijH914b8E2lRKJ5jr+PNVZGiTn8fXLJOORu/sYTJN3
NbHHSSshMJSqnDZ7AFxiwQd+Ho+5g3We1ZbTxDmwu0X6HMB2x8VOANXkgR+gLExu1e5BGobqzPf+
P0fapdEzDfp7L2bBvTIQy9Hj0ctZ/YqbjVJ9s1sjXJ5d8HvkS9CngN/9VuvvezTtW5AC15oqTK52
KvOl9SVnCbCsNUak7VPBNeWIc2/9zGX67gCkHDoF8CWojnUSsRAwu9G8xS+THIn6c6mivDe5/S1c
4RJk0XdAqPtJHUsU02p7WxQexDLF0vc+bl+b8H+koo9oOqB78z31dqOtHtxQwFgpl1YANk/E8mTY
RJB5JUOrXfx+jrCaC7MRV0Yw6VZ+w/sn+S7gyHNafiPX8v96MWiPFHU6GOgpaBPD1kUES3uPFJJA
CZw6MN5ewpjNswMfiTK0stADHZmE1AYFfim9MuRcrKcYbzLR6uuJxuNHuU/9QNMvYPfnKE9fjXlw
G0/8pMhxQ965aKfOkb/Z0QauYGYXfMQApKz/N46oViMMIQFj5JgsxuXQgicUYWSswZUFwEUllWXR
Cy35V+yFE69HS9NktO/xo4nE1TfnSCvFVr4U/uk1fVgQHitKyrS+d4ytW2zPKaCAKmgpeay6VsV9
IZ27X6yLXtH/r3cgBhvyDnNIY9tCrEVAonmlKgxCxbibjjLEsxiTDzTz9+i6MfidAB7AOky9xFxZ
1j5iBiIspVYBtOZKIF2SswhBxktsXwPi/gZkfBWfx5wyy0qH+E1+Lzd5DRysbHhpsqNNSkgBTNQl
zuPIKbdRDyhMOwZ/Dd8NMbDhEXa7edjQF1IPEESUCc/gr5V00OVZjBjfP3UakC4ZXdBIUbRT31Nv
3f+ai+ARGIiyg5lzIrhUROaUoIjnuShW7V+jj7k2ucy0oH9hZp+YfpC5EOH4i9pNa+UptO1T7SdC
ERCEUFyBPJVcSfPlyZr7gE0WzL2c1r7c1BR/hVlm1Va9H4zYombW7jpyomGe5I5VxS/P481ewSqt
IuqNmTE/e2Kq1X3TfgYWyJI6nbWrdHscda/NBC0RpOJxmF+FNbpQCNrPCMO+56bfLVJ9oQi9kjfd
QuZRi1KhXP2FXuEAErSVnGK4OHTeDXkuuo+K7hwtXG8C2OdjXJbYu8R6wcXLJgOHRyI1sEzgpLFB
BMCz306N4qPRN9bzsOHlTu+tkk0GV8xmrppmnnrasyUtwUdKHrNZeI6Ag57+v4/WFy1MWENfkeSx
gU9hB45H7izCojVEB70RL7H5gTl1OX3mVPhA0r8bD0RzcHELWxSqU0z5Z3RFIex7fOswNVpHG7mb
AjzCSZHl6wkOmxPhOU/YWlOlf7NdSC+CZCgDb+3TRkl4QV4tFfZiLYMQarFTF60HfSkteBW01/x+
QOsxhJG+ncbyQFls3Gz7hpgvz+nhqFYI1h9pOd17i3zaEc+KT2x3wJCA6IshUUjiRMEiMk0PAVvf
CuegNtVjqGK4rliA1tS0J9yks59s8Lb7P/hXWXBaZXOcGCUZmul0Tq2YvaR4zDsy/95Y8osRj953
TV0vi/FAOt6IuyVdgv2ZTqSPGTTATI0rXgZ28zV+PhrkG0ML0gAM/LFitdO1Fh8vhhWXdU4JkVn4
U7A/thN5h82CuJzlDK5WesPL64VkwFQttFutyM0dDwubGWZZxHMJolcpeTleF7Dk4MjYlG0Lul9E
YycaNnuE/s06yKwWsleHP+42KWJLMKmVEfdOTRG9ka2b9iYSJCK0GYPbgIG1G+9HymwDkkf5FRpV
geciaf0Q2JR6E5qAAHa09+6Nk8SIoQPaHc/MvPrzo1M81EbGRmiSpjmCTM7w2a15fVbc1nsSYMEM
0z66B4v0LUVP91x1B0UiPSZ4FZ915TtqGQ+N2EYcm63iafPi4Y/GEA0D5EhcvkflBaz1SAC5XEIo
g5RsA8ewn/0G+Mw/yhUT0DBCybWnnl/iLrv26TwgTZpdFCAePh0rXezqJNGOFqtwVK9ky9JjLyN1
9pSxWrBbDQbVDHA9IILTAR2WZhphZnQFjIghhRpW/4mSSJG4h2UshnUk+Ga7Y66VMt2VvmcKniIn
YX/lHAr7+8lH2mAQ2+7HoQV3jiXKVRLBgr6T3HDSrErx7Jyxlb0JAcBv66EaqcnIjYhS2U/NEVW1
TQeZ2jIQ07eMt4p7d05NMRy+b9icrPjM4HBVloQ0uBOviJAkTrXRU9OyZE/xjpWlgB44mXakUaK7
cVBUmhRzyxAJQVdxKmYTd1ujW+8+YyKnZ13hbZgnZ0YveT6Ezu1nKtPk0zMfSty99llVxJJQ6uXZ
7n6lC8J0MI9LSvuovf9H2lPcgLx8IsWGtA9PDPMDI8XuyePnXmw60JEOz3VX8NNOrZzH0s35h2Cx
/zujLBwcLOhN4HP/wM3gWQUd9wY1tnF7nFEUhXWvuyOVvIisQRQVPCIEmqWiX2cH/J+KzWKAGQT9
lzztrXNXCtrTqUWM72n0bZ+0ld7xlutqfj1rJ1ZMNkbzQ3bRH5VA52DRicCJ/jdfWTc4eyGxo7Tt
H//qw2X6YA//8sGYbFD150NM3cXztvuXpOygld4/ZIkUzPljT3rSvPHaeZy8RiuC2GaZ+rvCTsy2
H9GVqyp4XHb9ZYgmB+/LzMlleApmXqKpOtwywxjC4V3W7VkysJK3xpfi+bTS+7YW/BjjSdIMY+6A
RVkSg4JnYRTOUfluStvRo1OQyKv+6VjoJpH70Oy3FhFclQCX6LvCv9BpgxD7GYq3XJ6sYYEr7ULz
6ASGYzTtPgW40Ti4GvA7tTckU4+8aTkwDhJdeWOMR2555WO+ChC/73DMWepx2E0TazYUOawygmQq
kzPP5lpYmD2gD+HBUQE15yMWT9qT7ie3tNkk83oMe5FpxNh7y9j6W7xpg+Ymb0fnSssTPZq0+a+U
Fc8lmDo5IbHU1Ut9M8GXS7tRTbkR17tPSX8ULeiMwomqnE9L1gcZFocpbrmdKorxbbd0+hascYUi
c3gKEhhzn/bPh0XyL8VlAcEBdFfYgxukZRgden8TDHVcMr6a+f3fqvLDSyozm2dKNXJu3e2kWTeQ
AU1WYAHSdcLFDnTb7c+s0UFPuqs4hjaZHRSIkmLmvMa9+2ESN21JEHQ0fclJ6LVV1k0RX6bYSjeH
knp3i1KJtOFJg0dFvE2rjd0MK+ggU2OX/9RHJuIqyXRAZCZXIxxWX7cT9swMIK5VW6k+Sshf7cvh
FvhB9EdxNgBo7Od1qQkPIdxe7gFEkOxn5KnnJ9FbdkVrbgU3EbkRXIzUAZ8R7Q0u7kXHxG/BFVc2
k3soFR6O3vSkAwhOdpUFeOExM1Jfx9ddSDQLqncT5fvqomW1pqWJt8Fbzs9dVou8BSLhPBF1IX0x
+V0UPq/Lf7u+WK5sftsTyN+Dc2O3y5mj+y4gTUhcAw/QSY3mLy/VpOVCqi/CeAemBOKcVKxJvVmO
8cNmuuFYTIgNS+QxLEo/25D8C5qdGj5C7c8XnjZhv92vT7sY+NYYgxkny99khrgcNwmuCQyj2r3R
YhmyPCiC/0cjA5x5xbk/yWVMAG6tnuyo/1hVJhIoa8HHrq0px6eEes6l4r7JmPPzS8Fztfyby30U
Avk2pzEZq4cvfnz5qe7lUbVITQRYg+8M3fuJKlW5I8hHnNiF715qxQHSdkaSocxt+Yd71B2Ciqv7
fE7Aqgx4lJAjYu5LDdemBHcVpaGdAqG4M6okI23DoMKib5cuufoxaRb8cH3JC70lHgb/+t7f+bOI
glmuYxwdlj7Kg8xkUyyESxb2W+RTkQgnrXgzKqpE0uM2rvWd3PllTfdFwnTlG2nPu29Wvbd8uzN1
NnbS4sa8hAvxyC1oQZ542wxXDvFFZTYqYar0LKjT2hk6gK62whZiMmSlmoWpV2zQKySV+6L9xMTJ
trRVPnh1Aj8MkZnsyuFhSgbYkl9rRTHObUQxeDmeXaUfkMuHTuRwp4wNsmU9TXpkI+lzBcnUtf0G
dt1kPcWiNS9rMjLmWQTJb6PWOzebMu2ieUUljgbTk6Qg1Rrqr91wCTCinSKKqxHtpesHYFe0i60o
zZEJyCC8cMzzKhmzvuxh0XS37yA+UgxYfRYkYG4BmIW+54FanEe74Y9KYN4c8sd0nV3Ux5Mx1TFw
95lqF/WFHs/wD4Jt4GI220GHX4OyrWNtomelb5losj8SapaZF5d0l9FN1O5qc1gCKO1CEmdnv1+Q
ccM4NI3baTR6+Yhl0fXL2FxKV9nW1WhbT/uFsW/r37P26neUoJFYKxIfijqhMwWu7K/v3Z3iooat
IdRmerdXkVNdOaeqGnUJetSBrjX8DA+Y4JXEpPbSHNL5rsCX6BspaFJwlZ6nv4tzkk7MZCaSUbW4
DTz6eOER09ODKHf3rlyrwMOuk4tVBHePKhGBxbcyUFSNMyr236Vp+eS+hTeE2bT8x4gHhhJUFf6u
aDYaI9zKcrPj/dY4dJ8MF9OyZDJkYxs/6QRtFP/HKvvLSer7K1tZmxI8UGp+KLnefoXNJW+Mu53l
++d9EkVNWDlr/C2TeNMSQVi0djTUM/D9h+ybMZKhnu7s8eJpIb0PcspBkKHOtVP74PX41ZJE85AF
kzvbJrxiQu8ysL9HB3BNcfEFW/Hot//Cpg/Rlc/ci909bRF1qYB3yw8+1wyJL56lf66/i74d1euh
0b7ZvINO0ZLi1PXTMyogPpQocQA+HqtMK3QmHrqoIbfetqqrv2RMw8JdpoG0TpL4xZbV8S1JiPtm
pa0c6lWyenBWro2+X8lc+Xek7zdd3Z44t/nY/if3WIX4o9TclSNIESe9YzVqzow5YFLRwi46o26/
Zdyci0dDbUwDaKoPH9JOmONf/0zNrSdGni7hozffwb6nOtGEjLqzcyG7EGrN71uDaSwlxZ6fbMCn
j9Xk62PbOqgs5kW1k/fDXkfzMNKRa5IVpgezlhmUnlwPOVtRmKYVwSI1uXi5Lzh/ND+/tR23lpRe
qQebc8LGp16zvXTeBFG1iJqxQeiQndoG/q87/3qINDwXzjuZtDwPgu6ruTuJmSwOQVjBIC+GFFai
v40jj86UoKJZ+liDGNmU7lEzznUdCPl2rOf0o7khXwsSyG11AA7z/MQ9NFsH880KuXZcz1/OLyNg
efC5j1mf3SHg8i+SrqEzFIrZCfOouVMdQwle86j9ipGhN+ZZTtGbdCJg7j/yEx25pMz+hs8U+3r4
kT0uWNIap42V1FlUmqSdYsa43Jx5lBWwvS/JODrdAvXrxWIlj5pQOirjBuwK5I30uzAtvwejpJym
Jc3TB43lIXHsYXUisTC7RmN68CjdQzH0Ksy79eS5o6be7orcZBTREiGPcinrw1IH+HKTIhWaujtm
kCGefi1T94y2uKc+bs1mx+aFZriHpPvBSmD/B/c4TL/ZcX+PnCjTn50YNgMeL6JFzhBNIVWaU6PX
z/2G0Ax8vgpHx/7kLh4qfHWgRxV8CdkUMmUnTLbVyWDWjdUCYsGkGSty4xzFD6DlIlKBlRBpFroe
ZlXJIFP/oeBI8aTq7IwQfM+8yCHwQ2bq8hVbDCMgrVLcmofz230dGstPMYTXIyn7lGwU69tQJZCT
kP1WA258oVrWnDeOHpqjImrMWe5jJrvS245AcsEreE2NcyI+LCwwoHa53zVqtRsg+SzYovpoKVCr
Gv0SOcWjbj50FeI+oKlxqcMm8ROQWnATa16esOTnXNke49xMADoS1AT1jTy+ThPWThlbIu9fiW8A
NsuzjmGNb1fFmjIlMKLLxf2albUYHs4g3ikEA+wA8WihkU1KjxNBR9zlCJ34cDijE4Cf6IK+XIHe
7BLsaHzSYL2fuPWHpAUGs6KU6X+pZGkGQaTPKyo4Uih3gm43w2mm+tnMPSpZFTywk45Ba7DtDuYV
sSC7HzsDy19T/xiShGiiDX6JHZwwhGxXVO2DRSQx6ZzH5ULe/EslptR6vbzxOpCgfpObSYSRg7Pm
m1EVRfwCgf7R66gmJNWY9dbHWWHvNXbsrnqFWS/3R3Kg/5FViEGu8MFUh0Q7bCj+S/gdwEDGZoJm
N0/J0aym5XcfTuvoJFWarP5gzgPzy82qIA1lDGfIbux2LCb4saSS62iDS13JJyQgOjn69AptD/uj
sN/zCE04uev+4DhSW1zuOLmJwV7J25jTTKQEH4bRYXZDD3WwCN2D5sdsbuV8dSsCeWBV6yxEmPo4
pjNCRFiBf6JZuDcvBmNio6m/Kh+hvfIomod7vqyY9OUg2aWSty7NyU9a5br25svhdyRbxoCfNuVW
D32hKNeUYPiNvqDkCNIHvkU5AqqivTkLmyLwAmlRFgtS/JEQrp2S+VM/5fR0JwLrIn3K9BYzwlmM
3Jliugl//XQVBFeLLlZSsEev5Vr54Zi2p9xf82fGy6B+qDf11SMqX/Mqp7ABSvDj2i1JoKGM/BXE
hfCy4DB7BxA0coD6hG1WdYBBdX2ATUu1/L7QRz7eUCXZH08hD6QN+P80940BAJmhTb4TbZpSVNRG
SDmT2TR8C9Cela04a3qtCP87mihR7v5ZjHKhmb2LTBL9dCY0bM8W3b1hkt6LYa2nqFrqvWvLtKiy
WqnMojECI4L/ROtHwaaMziwt06T10Cs6tM04jvQIfq4N8RvTXf7cuOvKqizmpLkK5Sfw/hjpst1v
8qNgpkp/LCerJP7zRkOVCyItQdZBZunl0vD1JFjna4tvtldqJwk++j+GIgKPVEqO07ilrhJ/o7JC
n1Vm2O1D7jH5M9m0VwslItYrbeW4F5OFBQVRj0N5znUQnT3aaowEFvP9XQx9ShbNK41nSROcojbT
H3fLff2SN/7i1o2/S6CrIGkLVPOudy3hrlrK0t+uXfu4D02Msrvc0G+V7RSZbq4erVjdZx0Jbh3G
wMdJm0T6IPa2WppRCyU87Bf1tDjxSnU6373k7rPtOSLyBi+VEFbffpPyG+INU58n2fZ0Jn9n6u8j
KGGA6Ex1rif2yhwqOPj73jQ8lsdk0Yzpu/P5Q6qrpi8K/orWMHuoSx3jowj/o/Zn4Sx7Q2CsKqJa
ACkZJsOl6gPi/4upecPoavNfi8z+whUajCtiqVdOC03bDC8pIbQM8QB0qTKvnMTWbPA9lRT7t26n
XAsr0tUv3nNtdPcvnmxss+6aHJ5C1qLMPLzjdg+XwS2/HSV8mv/kgnzczKU318MYZOff7msCT0Lu
aazUvE9arp/Mt5SPSCmWRfvXPovXTCPboGvPRXJRhI1nNUY9sgUS+6ijtkIiz7/oT+rCT7J9MHAE
I4BfTYPpZvSi9m0RNb/JgvwtSsAhVOg+k2tX/Pveg+CuoklKjFnoLYY5AHnPpyYpnGPKNM6P9ldw
bQUPT83YgB630vAe+W8LoD1kKmkGQMLeewZsZR9CutdBySsnqCiXz5bl1gYt47WkW5ocuK8ptDUE
YGP6tYMsOTkc4rf5PPiZ7Xf/v3lOqK0S9cmtrS+kWHeA3tgx5y01zZpc7+ctzxheRJ/6S17RTwsG
o1EaAjF+ouM/6icLBUe8XVMBmErdLvzLXqyw7WgZ857so9Gd/YCNuGxZzfosiEUdTGqsPH2xZU37
OznPm/v7ncKdX+E0mY6e0VZV+ZXPofvk3Y9fFob2zyM8vztT3iolQ01qf+Tt3tpsc0vopHVJOJKI
7rJ7E7AWuePHPR2x9FGPoPLF6wKfop+ZfSsbdm4iYR6lW9UtUuH0huTT/T9bWAs8gFmSB72znbJk
z5t7PyRhuwBId4Dpsvq3EfJK5GmjnODHWJb9deNaTE05Ngq0OGssVcRlwm778bR5t37dqvytcYfk
QNfb0vJkk+2dtDtc0ZV1UzE1ZZwp/7i8uq/GOQ/LdGKcMPNIsY9ZxBTm6O82I4eR9AHYG14G/mTg
pITeYDbudG/QqEB7LmSiGkJjpy/G++od9YHgclvaPA6ToxHyvoMrxX8GaNB0zn/cEnYx189aZ2If
nu0Swj13374oz+KAs7689iTstoXx5pmH3dIIKkxheqZxPAgSVi4CMALBUIRKfmdhmxJsU16eRZmB
l37Tc5mdlSEQJKVknToHY/mvCUOdauzXkeiq2r8elxNjXSXZTDIteRmw0NoHWJt27LAdkZ63hSnd
tQd/HGQVQPIx9MU2jYzwZHUMqAOyzUNtUx1FsevT0EJ8NRICByi2d/Lqc7mg9wkLZu3CH0E7GhKO
ZlK/Y7f3V28F/T/GJ8JlOZDsWnDxiqFkpJuuZu/AwnL+84WBgZ3h3wbyGDnGdLsZNUpss67GD2Cr
ORz9o8TRnsVOhptftMMo4KD4wZJnIIfQC3D5N8yuAcM5PTinghDgl6IAJRVYE53zM0rKNeQj9iBW
vG/Lx0DDA10gw9uSqnd438pqtZshskorGNEx7NvyuURZvmj6EoUF6cmC6NELk6Ww7fnAWJgu7rIG
2ZxYbWARV+nKc47fE7H2miZuPJvSnkK5qMR7a1OHLRzoykpuSwppwbbxjiH1UkGS0kwrsLjEPlfS
J4jx1oWKAHtszTxBBunEJvd7PIwCiSM6tsS31dvP34sCGodLnTkXrMzNx+v7o72xRON3j83XxNBE
R8VQGo3QQvFjA247Twkx1xPgddWxcmxhwYZ06rp0s1JxgYcSgQ2tgly0sUn2thaO5IgaCBkwmfLT
VuIwoSsLznWtsh8Ku0xCA2sgprj72KsxY1llnpnY18B0mxRsuYHbXpGAFr7X3qU5cWzhFN6naKOQ
48+4CAk+v9y4OL5k+En3+fOAkzzXspbtJxZwMJqv/tYXe6Acv/Of4PlACbvcR3xkqkcrnByGF/Jt
2z7yN+4hbv0Gw8JjKL3g4lr6bfErMCZPSuPLXN+6TYA+9mcR4spOCkJ5EHSTdNTD4Jjr0F0hcLjf
NoOdOKU9289kO/El9m6DY1rAEP+zvt/p/vsvgvWjs3nNggN8X2uqEoS7imRTAlbKM3Kb3ABurNrP
MSk/guERtbLWaLrHa5OcDyMVktsuWDY22CMXySuFIC/khxg6qhwtQ8kbIJeZH+WE98jNLirBLJmP
MhE/hTRfU+wcj8aAhM/UpMHDdYVKkE78WlOlAhoY7B8EhN5ZFD8tJw6ixmZ/4+QReB4NsAG3sals
TZ6bLLrQBBC8YRMdfTd2MSeDVtQJluxONAo8Ql7OtZfsqIpEM+H5HDHb0hQCV20XBJmIo/joELUG
DCAMyRxwRmNs9YU7kj1pL013MI12BALGbCH3exgz0FwScQL2eJkAlXzdILHhFPopAmdKz2DzOggl
fPrttxDCzlIMlRwyfqGGtKOsxtpE9VKhHEQfcxU/8YiTP3Pt5fK013hLORDLpx399xuc5MRxCgS0
CWSBWudBd17rXL0LCiV+vmfOqKxH1luAZTMhJ+ZT9gBJ5GWebaBcm9i08NQ8ZtZZXGBVy8z4Qkci
A4tkKUVBIPOhs4tuLzRNut5s3QMMpIkrJ0Wij1IfHvhgMwvaATq6f91cj8LnLqR7c43uA0aQg/+i
ecRWoSraxBGEq1/33cGbpfA3Z11yAW47pUzC5cQXfpm2rJJ3zR2eV/Z1tX9PFjnnUz5CXgcDoKP5
Y/8Ii2MgzGyL03ojx1NOokCjRXQQaP98hi4b7EgFTY7hslphNGzcE+HYoPQt/6VWy4WP1LtDqwgW
gWJWHHH6e8n6r4igHJjICDgWcLoZ8Z5MwDRWPhRN4TA2GtMb1U7eNg15a3PIffrYRWnYkiXPbTAj
sR0sBTjkOvav4KG69X+DtzR0/ssz7ctjLVzjUJmC3LpMec2Hz1XKgD589VVYV8NFInOzQ3RCi72q
5tCiIXnPkNlLnYzslq9fVmLqQqBBVvJwQEb4JFCx/6rAiTbOxudFXXT70XS4DPoNfpBv2rMauJIg
iLP+szsznOr1yPQkZOtMgCe3d6TGnhBkINMtFwfPakKmgeVMQWcwTlniW7uB5iKcQkbKuiHVFIq9
D9+yYN+FsDBGZQYEWIdSvTMKPbPpIL/fKI9w6rLAGjYFiUArNpu3HKevaME02aCxmPe6UMsnlV9N
LSJgnVEmjfkTGJ8ESKDDrnCkJh49Tj2P/TEpMrvHBqBrusnM3gl1avfP9gR/K5hHnDTTlF9voq7f
HSZLltm+y+de/mPG7yVXqqKn6kLHOIK7vj/LlkiXIArxDwV2PyL664nWEUheOU2vGxnwCPmfdOBk
uNrxImWPsg2jNnlyS8iJmd/pAjZzGJVdZxScemiENwE3jD2Q4X4MyIcqyuV060+WxP5ecud6ZG0T
WNXXMwJ+Y04xxin2w1YPuy3aYiAcf4n4xjqq3yvYwmkUvHEcdAvr1hw1uXpH9OeEgR7ScTQ2A9dZ
VPHLu396lv3i/0oAMATGW4q6msr5PmB17gKOC/YK1J3COVAtfJn3/8Jyfggl4yT4rYG5r6iQiNnK
WCkACHGco8n+dOU0HkTcvidn+MYtcE6XXtm0/d2VqQT+oEQIPUrQingjzVBwQzEhoQdHcSQf4hWf
9pTToXnU0vVZqmgqIBfVolBMQigzJqapdrdFzjVyLAMvgvER6au5lsqQuhsmA+E5peaGKYna5Ge0
dBez4JRCKRiiWCRL6r6FGoYAvTKRAL1/1KH2HQ3ZjSGNgUTbX58bUEWjFgqkY3bCXBCv65f51SJd
PT2JjsDRs6cqdIJAbE9LOMB7O4jfSnzjtghzkN09ZLsuuKjGO6nEQnYMVsuyiNywi9GAFXEhNiuW
2KChrzeHFQ9Bs5vPAI3+PWHFt4dCWViZYCzG3xKUsPlEl2qVgz9ozD9Knf0qbu7OMSjTKa0f9IHE
gQA6P+cHZJ8ks9BJuc2AVFaeOjMeCsf776xsB+DlNHfWwWLsw5+y0BZTrh/7AdYpKTbCkFWF8LE4
xiCYOVsCGF8uzRKS+AACBSDKyp8Kt15dbcp5XdFXfWsfkitpIfyriTK7jv8bEcJoiEQ8NhWfu+hL
YjC4WT4QxfEdys36e2rgNNhUSBNc3iw67mzjo/M9OZT4t8ZpFCQDVWAmShBk80c+l84/dmpKpADc
A60+DtXYH1BvFB2bY2yMoj+r0zO9D8uwod5gTm7+A1Y93mS/XgsejtUue9KFqgmiyjprhDZVNzpH
I0jlDL1SoI6cPi1WBwjZNHjrGE1HZQ+tKTbWFHr0FeMDPHowacoGHFPLW7flnGwRuAdSZKtDuF7w
2wd/zjuIUt9RDYJJTJrZLDBA9hpPCa4bTSE0hTc+o7yqig5peBOhzvwyLj9EwbVvoKRRjQeqF4Xt
AgHFqpMzlyIUGWD+z3gaEH3iAYODzpWMt9/dqK7mrBjpHcwh8KZO+Yi1hA7/b+KwVX1pMacza0hE
TwG42Ea4PZvXHUCtA96yYYYzg+gdRn/3w77Uba7JiUc9c6RTLgYY6xFLTrU8o5+DInmsjxsY97ek
G3kqo4zd2QhEKFIOGw/SyX/9OkVKb+uZ8g+WYQLtgOhTK/7xVVh2vh6CaAleVsRTdk60LTe43zm/
/OumI6Goa0wy7BMvA49nrFagVdmKYYv68DBEsbAHTNum/oqjDT5apGGiHz8ijS+DKgpFlS5HhPt9
TzgxtyCKR95hcyA5OCAHtZTlDavQ1yCswkk5/DXjoBe3HePFFtk0r89QJQ2XltlXUia/SuQlTXFi
nEQRGvBx4oGiS9sDQcH7cFaL+/Y+x/eYN89pvO1sFrGap+oKO3uZ829Hw/hknxBQ+ISNsqZMYRLz
yLTkIxovkGXp8cTS/7sbNXDhkI2ocEslvt81svzg3f+YHI+/Mh1YAeUV8f04L6ZHebS+48vZ1Dbw
czi4fz30G8SdwdIm3x9XvjyHUYkEgvGu8dq/ttttG+gdEgRNwcN5HQWMBcK6jcVAEuUR7sHhAReK
rwlgteGoNMtE5yfdgC7MBYloR0FdN19h+TXYvPpHCCFABk+adk47WQJ6eVb820xI9LI+mq40VybT
Q0X1kSScT2rHDPkKu2/dqoSkQW9l8Fd5BHTg5yHyT5kVUOG5WqjOnOy1tqfPQVr356qpZBd0WO4u
P1sPpAQih4gkcxqCmj40B4G3bazlS6YrLuNlSsZThGzBBTE5uVn8dWvbISk6H7dWjTGMxAO1w3oU
iMNlodVaCcbfYLkabq3ZOwnLEFlr1FmLg2OdaF0kXSk5RawsxJ4VbapXEXHooY+1RtYHPHXlXnHG
4PLCqCKbFsG2ypHj/lX9hPLw3jfq1MeCubc/pu6Z64uuqv/CCTkabl4xxj63iU3yBqrBhsgjPEKL
M0WiIkOkVrKkAuIVPrfhhErtKZhuxNgtEwOYSoqT5Wap97UgXV8uq6O+0qSIG8Pvy+5JukuXjefW
EETbENsNxqoOOrlCwJonDQRZ7YmZGFZXRXAFACZW6IjQE4B72TPHm1awFujj65iMTGFcZPIXW9sT
RB9j/pZNUOH6IbI4tAt4YpLYZJtvlAZa95wEOT83dIqpxSR4vAoTi3HGE6nYuSk4XlQbMMamWjZ1
WpbssHvcDahY4nXWfKAvFIk/vds3cpGGZTXU36joKvjjEdj3o0mHP/xhy0is2+S4+MJxjvOuZ0nN
8f3ZC5gwYeGVQ9UKJekWQu+JAOXjktkKgHF7CEoIWGSahgIT0kQXbMQ1zUgXEDanaQooU/fBM4JC
5Ef+HiwXRfN5VbJsZk6rTuiQAEbqF6vGUQWWc7hteWjrUsh7NaCoZD2Q2ehLUCffG8Dv54etexbC
QKREWC+CTE1rjsLGWUGt4CWV7S2kOcids0dHUS1/CCjqRUVMzgURFNJmYInAZVFTukRAb3Jo07h4
Si5iSPeQYbE8OBWpWMCZVSLyZ03/zStf59D1QOvOnjaFDty7Y/KxMeujLd2TI8fU84v4cL0+UOjB
ODuj1iTza7rBamhnli1+scYNJxgfv3qpGK2LPnLh5N1VcT2CSg3bgmogq/q4UHeint1D0oKdFY2e
+XiQC7hJ5QqwFhzZU/+7WfvkWbjOm9jmlt6ju00494K+WsLB6Q8fTJMBHPCLX/RxoZyFWfxi/3dl
XObLmH6z/jywAXDIMrPX5It7l2iKcD5v8+NsP/GSyYe9QE74H9GUxos9qoffdnbYwGu0bV4XaKsG
qiwYrT5uEGf1NwZiAHQbhQKWL8+VFmZJNwW9PsOubm3Vw7DcJOb6kgIjQksriGypq1nab6pgG4qr
hSMaFdWK1Qm77At9O83SRFagc5KrYWlUhzulzDND3oO+zaC8dzZEQisnGsUP0OXCwqZMbvx7Xbw9
7ap7NcxpEtWZhNuaX0vcKtX6hJXjlVXIFoU3sOidnA19kB2CSYvAOngx1ObFgdwjT/+8fGyJL1Y/
9nOMKcuPtjQ+ea4ce6qpO5Vsjv4GJ735yOTXxFOhlI3iVAk3nL38eKj1ykrIsu6+BOvXvPdE+fL2
6e/wAIkjxvpBdZrBGwWqTlqsF3YZ4SLID233EtOBYYFBNVUMl7tqg34apqFnxfvRnuxWUmbsDguD
ws76IasXlBTa0tZv20ixzR3VfsQPLrMirO8nJLs5sXkz2g/GHCloLAk5zHAPc1d2ewbOYOKLCXny
enuHD7czRH/9VkggttHnLaLR7d2hqr0mOtb+Tj1Gwn6DgaWz2jHx82a79cJT3AWQX+GCtxlQkJ3c
7lBq5prG4JG8sJ2jjlb+ievKs3/YxSNQtE6TTpu8dqfgYo32tPf1Hm0wEPbq3JRVYxQPxijTAysF
r7Qeevrz7aazhnpkmF/rIwy9jIyL8BGAx0pOVQsIE2rHeI0Y0DaE8XRW513hykmpAlEXkO+/GxDY
3UBtdA4GYsYDWkg3JtxcExTyNo04R6YQmbofowAATb6jcUHef4oRQ7DHj8jGFIQsZBl17oO6v21T
HRbQoEYJqh18aaUnur/ZAFqMD5Wgb4zUa+swooc6J4SwXcSVBrrkZ/C9m54tsRWD71OBnd84fRBE
6hmZExC8Ykc39uWMYbnmD/gwGd3EQBP9x8OQs1S1MnDBCf5yrckMvlCfukNHfVUDL3zlVlOOYwUt
NGQQS8Q4sFoAaOcRcPf5ZTxgMGhcjRR6c3rwLDZgw0lW5XBf36qnNuG76BBwcC/GLs0pd30NOw6h
g/WO1nHESIOqFCofukatgKtAJsFq7gkS6N4Ab9icbzr2v9gj3w6KEyyD2AyVkRo4NGdpfTZQLMF9
SjRQZujMSPFmB35lCWMBCKUdwhu5qxV1/qGtkzML3ljWmAbsfom4ydKZkjYZCSdohhuo6AH25/tq
JnRL/cs5dii53Th/smUmSnYqLkgpHr/nqB8Nz9zppaeMxnrhL2ZU8wKsmMRro+cz6muJ6bkiOynZ
1Nv8ZcM0QYgSdVMz/205lhRepYWvzAGgmeNubxLaHE2ibACKBp5wHf+G05ERGift0ZLjR+lKO5ur
NBkojtmCmhWcUoILFo641LsjhjghQIqxmwfxLTeVDyWgWRxuV557Ah9rbp8dv9Qzyr4Of8zdaqcA
uyyjnaihpE9nSbQWHq4ZW4ZCXmKsUSLicjWfnS61T8Enkly3dhNuleujGqxnTdRvF3MF4HHBlQMZ
DTSYl0KPvZRQHNgtUB+Yo26b6CfHhnaYNFk9YROEkRkDyKoAJVOGVAUh7TCFc9BglBYpIG2IEVNa
OZUZtfi0fzk4caYwH9fCPbTA4X1mzTc+2sRqPZEPxWLrn1GkPIcteAdzkZi0zquSg+EOhOZ0Bzu8
DHa0IgzOkq6YtWxqzWpYfn3laCKVNbNDTNq/tZCIGh9vAfsAKIRsobZtGZs+IbQpJVlzBa620mLt
kOVBHFonL4xrEaQeKAqq+mbFks3nk2Flq+doeV6H35VPt5eM686xWrIJaHxmk04Z6e0OzUqdM0Mx
U1LWmVBMRxgpMIKUs/Xq9VSxzm+G+5pnI3xD9J6HIgGcqZK4VGC+aDOA0UQ+W/Q9IpsX8ntpDDXb
yqsG7knJGsJJOtwFyvHofKj6FEo8hp9XUII99SlGd1BHoGPlOz62FeK+M/4RQ9d+ReZIQoTH0pS0
OrNnwcblJUA8JbzmVgl/CtmvDskBtIxXcQwM0tKkIx3y5VnatTvRAzFnqPjcGYO4GIap5WxUWxIk
VGVJhB8ZO0Mx3jSFoimGN6oNHj1OfP3cE2b/PBsDd+L6iqMNpGa3a2bcGmDPuEXwXSxSu59qYfAV
6N8WbTHuaOcFScTUN+QRUJQ0oXIbl4SrIm7TC0e/IoV7/3HHOAwrhYCxEkYofAFCUdSUHWD5Hygz
jG3hoKX8/OR/o63SpbWO10XZvzuycafsdcpYFhZSiDsFJ4DQYi41sP4e8DRfgwcrLsYH44/9ONkT
2uGDaGw7jMuMY1UvjzJxuH4x0IZReqCqpQZh05AU640orHZ2wGWIg4o88CgiFm1CLHOAoJv8mIPT
CYOo3b5UadCYlK908r8aAl6exWakZo10nK59JesZP+HKoy8CIvVgwDXM2ayZ/ul6Cy7jZDughvL/
3lJIBdaFAMkl+xDPVKFot8btYKYMUrq7GX2HbP8Yev1JVmtQFik9VfYlO9/A0blwHDMT1kHfcXr7
FCb+3iRS5VhQK7L2dQjF3AX8hx5uFynqMJs70W1a8PEaYXfBalzhxedaHWN3i19BXOWPrWeGOWwq
YJqgsQlxKw+3qn/RsTgnUWPwb3voYGLtfG/jSj3piTvR60qqyZC0Y9AQCT2CdrU0ugHtQw+UwMdE
M4ipIIm7I56orec5CyFywJEC1RF8iy4M2APfUHSyq8evGD462OMJQQSJh/x20l+1+5H9By3xTPFS
KpjDylv9hBBv1Rs0tJQb/4K5r+yh4TeBy+LTnJo0N8G2DPTDUVj7yI+/d1/allIEYBCrXg78/ICx
/BiBvHK5yVV/d7dbN1kyIy8tx8gBkhdCqrcs0NISVuoV4kJEc7JOqF/3JMX551cB1knuJ5a0NCwv
DAPMwl5KmH0+mqd9w7KNAflHMyzjZ8YMFjHWyFF1AzNAH4+71T3UY9Gke8A0rPaTwj9MDaBd9srT
P0aZEvKFrOs00GmgtYIIk9cBb2lV+UD+PLtghe8kYWijUhYeF8UQrxpMD4/fp3UdYdT92Qmxzwru
qwB8FJwRKWB/llbdsfn+vAyjrJcUL2Vnq9+ZhPIKQxXK4cubyffioYfkkc7cueYNlFR3i/uPfXKD
XQR3pHq/AFzsIOWjvgjIEX4mr6CIWzlL4caJC+/B5Co/POaXbuEKIyE7wi3ul/wrMoyvgfau86cP
hVRTBSffuE1WLBZQWCPAhEZCHf3SlcA5upm0AkRtyTVlVczoi3tcCCxmjh1lQpLLg6EBge2C9aTj
/Lxw/n0Xhs20cU/I1Ag1m+++MvXK6HJKowxvKFoOkf3xcqKC85vmvC1zC6UGxr4vRBOgRX+89bWG
ya/px2OsXitJu0qEk0UbTzVQrJG+uAZJ4gIfB8hBObxtuZyUuTdlgW9hv9hMbj5C13uzq9agTWVG
f1RBY+1/VWRlbolShMRSgq0MpYgJVdOFMVELcF2rs46itXp4vFQ9LbaZoV5nDKPQUYJkNpVrw7p7
1pJxk21gp9TtDgMKaD/Im8l62DCn8mxXkL+49fOMNGIEo8PDemW6S2tmuIYRieucEne7bsLq6DuC
6ili/jE7YLkMGNvP1OTwREf3ZGnd+AFbpYchZquN6S34Ob9GheoC7KUeWO1pX/05TysPRKjzuenP
eA6vrIzVeYexzBkcNdfn8GHCqPklgzOfVREpWB60GY4ZEgyIrmCM3s5AYIZYZ3BKE+Zah3hCrYMq
FMph8tcuG/To0lE822kpxwgvjJdv7on6jPSrAjYHs7A0E3XkC4JX14GRjeHHkMy12C/knykhVw9Y
2JzwCzMhs0znWX/yY0D8tVrxof4ZA2Y+6UoCpgq5g0I6cMVAeXQNLs/EDqoXM8pnJTOhYO35yH8m
27TCdtg+tV3QZLrw6pWAVOQ4b1fMNLXajQ4InEAHSOcLSafeQZO0B4SZgpDPuTh3nvIIYkwKSZd+
N77Ha0/zubb3V7K7bg5iZMfiKkVsJ8M3H4UvF3qyrSXpNjmNuOgx9CVohDXc04NAmHOO9NCcyUx3
FftZRvTXx4nwwu5qA69ZSyT//rH4p0bNZkRSXgZAAYJ/wn9MH37bc7cbc49yXQ7g8eFxT8IA8NPL
KwQ9ZhL8K30iGDQfGUk1IeuGyk9x+mAEeLP5tpr437i+qaSl9ON8YrxnirtnInX/GTtv+iGfcrQb
DeFVLf2da7J1p/xzlgV4Zl6a/UJwJ8B37X0NIzYJFx9U2aR+KAS8YZITSkHLWaZviIG3+GjKPC/P
TcnED1y6NtwZqAv8hk5Z/K/XyjkvmaIdTMNOWGUG7fHU/HZESTajEsOlphTyAs4kwAsWTdJMy9sv
Ymt8xGVNQODV6QqwVMft3km0hIcovzTpmlwfSg3YUAwbm6g6gfUWkXL90Dzrt1DanOOvT1xq/CaR
1MhqZJZceObnoCOZFWPhHDm/JNaxs8dIPlEFKTHjYRRfGo+RH3v0osUk/noG2FYTkrVliQxFqYry
QwweWDtxUmFc4XHo/z3s+mVkzyqepzJZ6jnCi7Ak30YUu+ra1W5Euvb+oyl00Bf609zXZE4Dajgt
YieQPwXCj2I2EmdE1H+8k43TkWYUq5ZvcGn0ATfCkbvBZBzM/ShP4Aqk7F+XwzwTyKLsLkG4GCw7
zNkkIZuIKj6AJOM/T23SoB/GeREh01BbJj1wqvLGwrcn/+TMNDgd1i4/Pj8MOPilZw/e9Ojy1tCV
OQTxZaIYw1IwILnMzODX/E78lod83YNyHuQUtsey20Rz4oAsJbYmoaWoUlxxx2Z8Xcm27AChppAX
q3tm57o4mie5JuqXyhmr92PqlW58ZDsPdJiIrk6FniLEw0dhd53hKgUtRnhTE+iRCNVo22apzSBE
vjGyVMk5noIKNKRKmhTZGM8VfdrlSsS5/yNEF0RO5UFkMGxOl80CrGXLI6BZ5jwh5ZfUHQ40wF6e
hxjDCh+NKoi/iIyc8ScU5LuM1SsD9kItKycTP7erY9OgdOdKBaIJvSMgxX4JXC2x8k8RK5UAXT/j
gGwVvDdkMSA6bz2wOPnSViDSkPZjyzLbZRfBA5S/aK40ZQVTyHfPCyrolO9ZDQzgScpBi7rDgTLB
5Bg6ChZpsziNIzZwQtQka0XW+FHpWxfrpl2iT0D2Dfcljea0+AJ4FxZpkH1Jp5i3Ol0SV3j29KgX
Y1DuvOPSU6e5pbrHTmkdQkbGoPeDfsGW6obkuFQMOZZLb3mEJrdhxffGBeI7LDZFeR6YtSO27OQt
NJ+FBnvvI/jnQmZXvz4UTuKKEW5UEbcIVjYrNFmK9lQwRvr6pJQYiprU8nuQRZdeLagVT8lzoReV
udcgUAeiVAMC/NPqwzRaCWGZjK3MRowmMfiHsZLn6967o1zG5tkOZ4ZmZVv28ZuaJI+Nvxdfdi88
zkj+Tj7MFtvG7rP5f+NgnXvBCElJun669ccL2nelxdoX6Yab9b1bmbH9Bah/2gvrEbGRWtuquz0k
yrkQmom9PG6MoDs3k/pa5dqb4cd7LB8JI3nuDgA2VF5KIq1Yexm3lvYcmVPVyI+WYdXaUsICzpeY
qG6cP7pc8hsCa7WrAvbmTtKhsxVIF/b5N6P9w9Nizs5eP1BYSiBH1PPXqY8iqY2QcgVMHtOomK65
okV3NSlYm5ncPgwRhCx24EMgi6PEAd+lg0sMXycilwOiHsGUUQjo8h91mifh2rsKOgTfN54vaq5b
BNyJx0m+nX59km/yXogSI/LOyTT+HG4+lydTEUyrywlzrKnWUlsS86djb8GC3P/4pGVoGp6GSaCz
NiybRDBM6dsBcvXbV0YuG37n6q34cYu1cYT6XOtnhISUu/o3isTuUiAuLWMVKVRHtUUYjRL/pF2B
P4MaU+BhIhAlfClYD83hW96NTkGA8ZGmV9op7C2dzNWWZ+FsQIlVCrNwLbgO13hdlBpC1bW1fRI8
5/AWPlqxIJAEOWxFAz4bM68WYr2rpa0fOkru6BLbVKoBR/mpWjEQ9z0scIx5skeS5s7v0/CIZlZV
sklwZlTCr7zFdnGboebXsw31tOUT+vTeKY7z4r7oAiVoTS/9ouH5ePQOgjXzYy6VAJ995MB/LRIY
0kooaAICK9ka/MFM1x1FePkhpZqb/VNCEky7IGMJwySWol49qPOOM9I5QkT/HvbDy3uxrQAEKQuE
rjBCSAQLoo81VE/0fPiokuO9ne1huh5NQnoULhpiMbEvcfKE9Wb+16kSxhk/mv9h1eT0LyppGHM/
OimUtavGaNDiZRAeuMoH6jQkBz00WDUvJsV40S+b3HNlCI5h17S8AOiblj8li0lj0xkbll9wxRmP
rJvw2UlRre/H1i4i5wDrLEMKYdN59FvqNI2FcRMUfSQdBf8SYXg4gfy/gM9qareRInA06jGKdhv7
j1fmP9oThSA5t9RpNpfdHZ/IMn7ZRW/YAC2RkFbOGP16CWN61I3LRbIRWyCB9CmleJPoU1emuV7B
f1Y5D9MFyafidZn4xnCIUfjSJg9jY3Ac9pkM4nYlH7/x8XxXEbeCxHvW/0JDYz2HL6MtpjPuQrRk
XJwxOp6e/goouI+CNS/Fsb7fO4f+NEemiEd8W92nXP7T1dbyWvXe5BNQXglD32GbMwgjgB+n8TyX
DKCmf1cmV1rMyDxibjbcZl3qNKxuY0CPxDxKrJ7jRdNFYYzkYOKJVAgeyEBXvL89RFYwjzZBMaZ/
A0hwIZ4L/RRu10RnKfrpTLbJqZe5UQywV/1IrWVUrLRyIgh9YuySmu+l4VCMqhD2+jnVwo6cvyES
RWFk8B0+CWFBL9nmuxrolYIGvvYJX7evEbuwV8AOlAFRt2W9clz28Qvd5UgtrEYQhZbYDziQ9ei3
L0AjQpmxwdGFzCAMW/N3gZdSA7PIgJ6ELH9Vsxo0P2Z3GQtB8d3RUNa4YKdUKvij0qafXwIXbbVA
P0APBIwHNr5OAhRtRwxeM5+9JRgHTBBEpmCgi4tf0iuPx4NUUvSOAmyL7W23UjQpoSCcCeCmh4gQ
mbc28191J1HFlko/7cejjKOaFwNpPOoGLwzf/aJTmhjZFH++Sk+RLTycxxnKAfqgelVAg+Cl4APM
MoHYn1T4sqy1tUXS4ZpwRUFcI7tZFifhvJQ530xbGt5DIlkFwWJ8cBTPpuNxhle+4Tw4kidsjiNJ
CyBVIZBsSg9/hY2xXNznsIkJGVU8LTvyBHky1cuf69nnCHWHfVQhyDd7x3r3Hs9aSCEPynk/oFSs
uN5fiikXoMZQwtXfp/96WcU9POKoG+SYRFWmMCbligE/NlqDnJlGgQWswPA0Za3vUBM8CzWFZaG5
M5fgXWF3yLjMGOPwXSyhu3w5EnYPridnePYP62bOg7R4AsXw6bsJthX45uPXnhPpFOhrWrezOGWZ
GYloHgzbWQyViM0XoLEsbO5WAO42lKwVx5FGavTUZabD2XZNuRHbMdXmrAUe0Hrd3EUvcIyG8rBs
mLE7VHisYA0HVHyov6cUsPXq90YCf5dMh2gb24oTIQgBkNvf5JqrnqHbFYzEf4mbcBLjtdorw3r7
214NVEr08YX4Oa3vMEa3/cXajF31iGH33mT0JAOf6LXb5/kAmjXxpHcGnHXnE8PQO6L9X/7hmIZK
KgA/J9RN+PAsokF8UGKZmMQSYQ7bor0n5GYy3AU56OwT2TaokSLdDhadzJGYvjZTbj6NvMEbKJwS
ilXG/HakdiLPugz1upn5DXU6cq96++UnNGvToUdXdihcvzVVvVxIsSD7MYD3lIA3kEu4ZVdEvMq4
DI0X7B6ijEkw61BeAleHW76SIZH9aT9OfYjh8oRPEJHK5J8aYguqlcRY01uOcoxaM80ORJSyH6Ig
B/kRF7kwvp2fAxaonajTDlpLxbe7Rc0akUoDgWPD9D++vQF1SidGMPHajlgZo0zcEyRNjbe6pg9Q
GGWpdDVxnQ/AkiCrWxV3Yk8owv8r+zO3lMK343a53uqRcO9HFEGuBXR4Jt3iyk26bAqVmxSGNkjv
yX2gYSnFRWzXrDvwwPBqQ/k+mPQ6UvvOLaBoPlqpnwtRTBotfNDW9RrCaedTLLEb1qszskxKqU5M
xXWoHme1bPPrCPUm+Q1oGCmiAqhrC1WSQ2+NpSMx5Zg8wjxZlifkHmR86CReGvqyaMwopuBhHsrL
2YmCK8zcoYU6wNz7Xf4wRTKrC4dDpFBDiqfR1/D1xtRgIyWlGKEoEJNiP3t0XtoMheqkw+Qr4TUE
vqo0RiImCQ2a+RpoI0BLWEQdE1JWesPiFcRX4voqQRA1JoUibEMSCjUs4gmptFxLhPWwYfzS3hSW
3FvtuoVNZIduJLuUADswJ6uVQ8+eFxj+ulwr2AjBWOvZh0syEmvAJaUnnnDLNKBKSJOzlgOfRBbw
/qT7DXupMP82gLm2kwRlb9AFf48kOpxkJqs7A6679/B3HjSvfEkD+8S276TH3ioCKBSdZlrvYyQ4
7Aj7H3VH6rnGwudC0cZosOCGa+pNPjN82tZZb1OOYczvSMZH9R1Z30FVRhol65okGXhV2AmxN2tC
0nJRm9BkU7rmRmMgzxJLzM9g/vxsBhGpbZCS80VLh+b0rC85D70jeJbX3XIZehWfV9oAbg4mii83
Jua0rHYp1dJla7GZkL+RHPMknxvLwA2zKmlyZdNw/AThkc6JUkYxcgKm4GkwTWmsxkQ3y/8iVeiv
NMlyQ/vMD5R8y+ynG1030NvF8GWxVX/a4LWlAxuWB4V6y1DgoGZi5zdTuWNR9CNfZp+geq7gaw8B
ep7LDTawG3N44Pwg57YzqNhCiNnMhSqDAP2nybGLefEWJeSj+lPLepgZ15piOwGxvH4lv95WjhZY
v+xDJV7ZvCa50p7aLugaGJO5E4z6YdtS74BmMRN1Vx1HsS7qckJbltp/34gHUT/8Yx0Ay0vhKsEz
bwyZVrCwxfdn27cpyy+xil3xpjjuQES128JBjQXblXsMzSBiAHXyfuuTJ/0xTtEAJgWM/998gBxo
cP0MMnzOAkiOqrgearqjtxc8apqAYfiGopGcA4PzvyHOp7d5l3qr6xCr1+qCbA0hPBrTf8rUhTBK
5ZQojZ9NFlQTulHQelkfAP+qO2+NoHDAoO/yCHeysWACYTAhlZUrlOD2g3EUY40T3H1a37GBQAYk
VEkO5GWuIZEyl2lKXNzBvP818vt0pfwISpgLAy2AxDeFh+kW8FNxxf+QtzGkRDeJivOgFLf9JRoT
k+9Yo0Uz3+llV14mEoLjBPKyfak+j7lI45tS2llx3fM9asIAyXvDjGTKm1Bt48QgPUpALOIKkzQ4
/yDFy4KX1iXuv7rqZytaopvqCgmaThm31qTZCNoUCqWPIENPiB4xDwpg8ucxeGmUI1Ft4QAQRtE4
w5ycj90n8tjZ0gq9u1qbHSbiT+zX0Fhw1TIjOauuuNw+LckThGBvgG+4bo3KVmNgRwkaWaReTtl6
+IdtS7PHMyUZZpiBOk/c/ZJ9vq1PD7DPbignYuPlvow4XgODufAzL7to8VBKrYhI4iZsz3piblDb
oUDgebR12d7NR8PnrZ9fwgTRZQD/zBW3wfghHxv71UhK9s74WySHjgH9JytuimpuRoVra+N+uQYr
0pydDAkYF5p5kWcrv2tiqsn55Ela8CtY5zuVYKLpj8hl0S+2z3Xg5J6XoM9R4ukn2NLmUOumZVkh
geW23eOavRH2XsEXMv6gkwx8efkIGeaLQu5W2BttXwOrOyDVeo3qRyAmYD8wGJsRgFysc0LIeC+H
MUdjLp0H54JKM6WXWyxDD40gtatwaGOZvPiA6U5APCiqGKVkjpJOkc5KSKY3hLzl1xPEezt8B/W8
7RwJ0WmMWxCPMY2d96VEaCJGtzlpf3AXyZMZhgxGiaTSz804d1Wg24XF6jBQjQeWgL5NHte+2/j5
Hv3P0lD8YSJPT4mG0kMP9llfprH7DboRbJEEmw2IlF9s5RJpcE866uumZBigfyzEtZjUD6GVTd9O
kWPzK2+4WBygeT+637FOoEorzTNFwpostZM9X/JZalxz6yXLo5FCZ9jfkRxQScZSRwNNZ11g9tca
nd89qUGNiq1arwn+Tp4Xi/1UPVKiVuzkcAyThqnklquLhsq4NwrrIO4+BOc05BmY+FzCbCUZz838
kIlbic98jzetUhmlwjsOI111cBXHQ89hMS1y1Z0L1Yr6MZBwyZx9YahZ826v1dP/tm1nhzFXZ5Fk
x7Lo7Bxxg4WFfwamTHpDVrZ4t8icwUMV6cDGfxMEZnz7ECgdR+jr0zjLCUdg8uGSqbR8x5o+Z/Dt
CpJQKWk48we2rmQnCITSuIPW6AbYOfuSYTDde76O3EdOw+frYK2HRZWnkflMJQkcyFVsnR9IkgFd
pkH8tAKsrZZjT8a8zv8Hg7GB2ER0/UBqL5DA/0IStbNj4NjgJDlDi+U+U6zycvn8FTCHhwcrjGsb
H8TabV1pyCzYop10+eBEtRwtmUN/zh7duA2k/Y1MvtCJLoOf2kQq8siHu1XMuJnzeQc2KlZ0kMkX
BU/6UuNMFfJYcYNzqMzBmuAklR8id7D2TvlShBc27QGYu5q5GoYUqcCqkjdwQOt8Rasb4moyPmVg
JooJzSvC/R9iydoNXPRNmIHToWXN8hGSslNd19vM8SbJ44+QjPRwT4NZnccD9Rr6sHUPEpfk2PtN
Qk27vlVmBvSllGQ1ZUKQhkeQYhP5FEbSWB31IubD3Bne1m+luB0sTHXibH8JDZXwbLwRRxmEz9s0
u2hthGoETkpHUHsrHnnCvkUeD6a+QeBh2mSTAh/bqCd7aiVx/lQ0bemRFBpqzH4m/ydrWcEM+40i
+7/Q/B6Of1ysF6JNas2xr6NGajRn+ncmSBDkR+5hPNOwSY7p6xnfqCyaqbTxNJk1JzqUM34ofM1t
LLehCepybIINajFDkDI1oRMv/al1WZ2Kl1TGvlwtvOr1ARkKJw1tuVw524H5dl9f6eMrKdwiAXTE
NB7lsGKeRQOpDoXiUzVknoqtQ5kRHYnrbdcCUM7Nq8HINd17c1f/LeVBrLraBQ7Et8HNHmb5+pP3
KkjwYOzoYSgqTPtzsVOXIjpDBnETE2Xq6Kq9XPCgKPiR/VRzxULdVs1fYHvur7YAqa1/XfmmslKq
fv0YaTTflZyxSy1a/tN23dO5LJG1OWwQUAb0BPQWUs3KCvwN7OvRMyuLwjyb+/QQSTDjb9Nar0wl
kxz+I/v22dfysStRC5dEQnqLwDOIjli4wF/TZYM/OPcCpNN9S2LoDR45itd7OwsS5qFiIYUeQvC6
KbvLcW2O0/zGGOMioWlWChfT3XvTHEtflUrekL63Un7hkPGMjBRGgGCWG8d8/tt4K27uCf5pPn0q
bYqMn39CIyQaoU2TMjA2EVzPBuJ3Y/y3XBH2IF078Q8hlER39sOR7c3t8akEDHXaeSHFyEICCAcp
aRJrcsvhJUGUYdkfHuzCoVnlhbm6EQa2Q0SZs7RxmNEeFk40szzPoxtZMUBoIVcrcoF30Cj4e7kS
AJBdTWzUDXGF50j6FLYvvHI4EfgMx6kIgORwwxF1XSv6bHohSkvfNt0bwxjhsi4+XxsTsVc2YPT2
8PC7g2iEmn3KYja9C1d4AmctVlzmZeLk9kUN8YJhj2fwxXG7c9+yE3I/3ugd97lwPL3tw5j3XoAc
z1CYdPfMheSKwRVm7Ef3G7o4XxL6ok+ARShRWtO0P+2Kyxme44FiNytaRhB0UOrG3SN8IX0UFNYR
/TL3yW+Hd7nl70UU59tWF8bFF2foxVes3v9yMavyWAV+ZzoyF38sJlZwRdw2UsqNYwSTlKgaTyH1
Ebf14x3JeDfJbDi5Zs0XRmex/oOUb0djbgST7K4ufo7jeglzWpVmoPgnZuXNiTIUwl4NbsY+vsnk
/0Rs+pZexNtpu7N8getPMn5jrBVUjIJT1MD5G/jFbaX+r0UGoXGnv51FC3J8P0BE75PEUuTFwt2j
fyOtYyFKKH7TEPCqB5li77JefCxmXrJ9dI5joJqMeuU4WF5uqgyWx/549NZpon9Q2F4bUC27o9si
ilHaahwa73CJBO9rVDgLoKWl7KTEIWOynpTD2wFeRnOL/6I5x8iNT+BgFmNDEhOau09CRtjljd1Q
HfKMlntCtTEpoFnSGcuDGlt0SH1CtNgtztuAV4tf+0S69z6GL7DcpuphiPQ0aS/qHbm37CSRsqQP
wPQ0KwtMMXRocQySCdAo25Ay/xegy8gTmoswA0fuA0JacExFWmfMyqlPYGjeLyqYKCXUrHzlHGjE
n1ZToYtD4U0UGVkPTJhkAzG0P6kmh9l/lw5mZ/MQnZ3zknioE1jwieRz3sJpcuEjnl5xgmrQC08J
dEXhRuOxOdt1LNlQ68jY5uJ1VsfTHOm41eFY8I+Uoc9Wp9NtrrdW3H53ra79/PtaIycFi2awr0YI
sVOawnEYKICu2cqULL/i3k2jvGhvW9CrNm9Gs9SW8K+HTpY/DdUFW6RDDw1qL4rzUXrVrFRP7K97
skrUkRum05M10MPfQXmjwpqobIPyOBxBaAe0IVYIfs4wobjB0RDWMf5EAkh5f0UmIQNngGA4QtAG
99LALe0/A59oZkxHn6uJ/HUP8ITezWNq9YYe58DPWVNfGZtwf0nUUTyquwidjSNMKHUKQGg7XEbZ
cFLoeXOHNuqGbN8QiTbPvxD4mNvvvXEA4TJaHiEMMTDxT0xhE7xKQ3QRnf2QGkT5J0QWlV0AqE5z
ImbgAeDLvvCU7vlvAhCTt1y4jFODGqMx7pgmpcpaPda0PMRHVACnP5aUtWXNESE1HyLbwlpNXEyn
oZrEU+4QxGTfphUJv3/yTGft/dKrs0RFm407ZBMPoKMhICLETZDqWhSM7oNnej9IzM/NWbCzDZ6u
tjQl+0qom0hU/kPq+CoIuAhiJrQMt9KGGX+d6dGn73/rutNa4g6qJIruM+gooNCZFHf836jc95Eh
v8iFPxxC2jI38ZbQ9Do5Q4BxQ3P6PiR8039a/BBr9c8F3D6/GNBp38mm4n2f983XJS3cp1i1oanJ
bsKsbjKCwYXDjCYFXsmc3nwFRoyTz/vAB4qeaJMOWDqsxw2mPe9+rQ4gtsML0+9fSxO8Wbf8enC1
xP4G2Kao95xAzFJkpdHP6p53a6eC1dWUOuaWwJ/QGGYciH6nhtU0sSJ1DWkHm1GrgXbn9KMT5QBS
hmxbfYsjIwxkWFw9HZxJT0HwD3w5X2Bk076m2smUqA64Y+pYWVIpRx3UDvMcgay2sF91t/ELzF4w
HlxQpi0eOaEAgqKDAbgfc13oVjNBaCPebKOKhFm/yyssfB/Yub9m9hfIV0/bO2kqI5Mdvo1izhoa
Kj8Pbala5Y9o8uoEdtENeVd1dcA3cU9qIl1lhPPqoTLTtxpsarpaPwIyRbS4Smqt4jXciJ+E4p3o
JB0waDsVTumf2AcjjAtzj7E40SXiH/9av6Ep8llqg1klYxOSqifB3tBQZmeBEnF2vhqLNihzA5Yj
gQVis3vU508OnxPI6iJVABjgcKeaKtY1wHy68A7Ec6GoV1gN7BamSLs3QzFR0TEvdH8gJ5+IoDfb
3fjsHKuWxBqH/YLi7r0RrBGCX5jWzDR6ULeGelmLTq2PCBTatXqprEVeLVv+L/3e/hMQHUbDGZXT
X6X8k5jz51ZvU7eF+voITG3tKSc/kJCsRka7lEKLuBwQPq44NRTLym9jaAbg4B+Khz5LnSz7cYsi
i59r2xBHGowNEcOKpkuFQn5mJKo/kNqMV6z+E/3EA+xDyUOe1CQmDsxo9g8uF+PJjG5nft9e5ApY
VCmJlO9qXudGIX6vcPApQ4Lfa6mGqO+ZfH+bILoRsfPEEQ93D64rcGMSTOawW/xRXggbFKLha7bD
/BoZX6jAyZQSbkmRunXYsLFuWIYG397BeYE01YGE8NRQNiwbfyaFBDbTqCuPgfxQ8ZPOr3WrnDnm
laJ2rDNQVKJF0mhiVrKzuuOm2QXQr3gqrsl1VB79APrF0pCuEBbqnbN/2da3Swc31rLMJxsHLeDR
jt0UliS2dbPrAbYWxy9gGSCTzynHUgGNp62sz7o3/VCLSCgd7Uu+hibx++U3jK17UlAPN0vmwW5R
7XJ5FiGTStdtx0Z9B5stjuTr+yH16Td9FUVQnISDh5LogSMAoQxFQzWQPXKGv/4cwFngw1wDPJz+
dgHQsXN0aU6DGNr7lKiKo0th3yu40HENaGmTNt9eqh9uBDjGeafK5DTOsl2VrHKYrww0hRDSk99I
lzmIsH1ZgvJCmrWMjAaiO7CAE+RPH7VbjqmrVeyjKKBcFIDKdUJMb+XgMLyYeSZRgpl/UaTwYuse
AhTcfXR7Py9JkgkpjjkA9DjQRQ5V6oY9LARIX/6ImvvC4btxN4bCRAw19X7MBThCvBW69F2udxex
ecCuRxgqqY9hM22VVtD+UE4aGM7IvLYZl4rq4697Mz3c7sym53gvTEWGYEHs1k1EdejeyOlXp/L+
8Scb6VS4YJE5c9D4BkBgImuvgnUyV4knRPlBfmSNCJZIVi3zQUO6Lna1o3+dTWwiB8e+5GQizcMA
A0s0dAUa0VvpATbbHE35RRy+3yxm7XOMeQxPCCDH2WcGjQhkzUE4rTUEnXGPeYbDe7bkIHVEbTpq
reaPfvGxklwnYSikFsU4y9BENle0/1Ma739IrJXaUF8wakBMzCp0ZoerDnjcEyIfJgdYzQBg8J6Q
4QHZBKczw+olErAI+nDkDH+xK257OTBQkJH6/LdlCL449oKdydpuHUIy+mhJndzpvrEkxnpCrh91
CcXBfn3jvxHtd6WXQCIT00kx02pz+C0Yo4N9oS/t0+hHJUYlhiH83JkP3+sn89F89cWqBsH0vDDs
dfAM1gwrT3xx2AMucQdpMsqaaUGTzImUsDowRL42FkLyVSSTWLVuHjpC1HYL3ioxJloZV+ZlqHsQ
j7XaxeuFxKN9BFvhYzS5GWftUOv2sf6XHAzWuMmNDge4KU6sGqtCTOqe6l/zV4xSG2TqgKJ5Ov11
vfpz/To9JAB1UqeS2QKCY39EmbGM0SPoUlhjXwCBB42zAcdIFEb2HQNNl6A/zNZmlDMd8IfpOKCh
9z1K9lR2UoxI53FTW+cgxS/2F4yu+Ds3heI9L3Ijb2Buj4rHr8LaKidFutPOPQmhEv9CyQnFCmfU
+pXjgS+aaJczI6lHH4gHdh5OCRGr6uRZM+tjo2hZc0gGgmpmDFFUlV5leAPnYktmYCd+1UR80uMa
sMMDg9IZV+dD78CSpGE5NSL1dBfktQ9k5m+DCkAHnZgmTTi1N70QekAZtAxC1g94GlQA+PXim9uq
xHoGjEBM5CFNGjX850HGzyP38+zZtji614XBJNXbhisw8On7XYgOCgRnE0gBjAvgAZhUgemx5Ce7
EUZngMyCR7WKK7eV7gj2sjh+0RGfdZmqKnCiBwDOe8MsDqkWuU5JUhtjKNdv8m/MQUpY6Fdix2wI
y3AJNT6ReNwkgaeIi/egdvfK+6GMlRq5K1LihnSawO2Q+SWTyvt0pR7wRodVR2VOIwDGq81/5ZZq
rcHAoIlm84CnheKNZSbGAvYMUTMignqE849NNmWsyraf5NJlxqRrms6b7FWtJV8rqItqkpV/Fb4M
e8Gm5OpcSDIArAi6HI0IINZWj1oeXZIEB24q4TDKxdq0/82+ag6GDLJuS3nfW+m/Bw2fZvxcQLKA
nMcIZFus40x/NgOLUu6dLq52W1QR/beMlUR301OUoCXswuTVAQD6qHhr0+6KWa3UqJnKnv6+LxSH
enUSlLaXsIYBPsn+Wo1z7ywrFfn15lYGidFmRr6d/ZS+P5WJL0LKKqvyCehnPIQQ663tzmBI+xOn
qGYpxPAK400nv9Ks5SM4HnNYVdSHo+a/JBP8iJFupY8mWGqgvTfjWjPZIiKwi+C06BPDFOOIdE06
iW813+6J2FLert4Vang42QjYEA+ex+tfeOG/zvxDwg76tMoStl7TMgOBJtHe4xYIlAXVCHRiK3H9
UbhA/99S7I2X2PvvQ1CjX4U1vdCquR4A9NDHOavoehGlRv2L0l2uMiOyOdXR/b0O4KVqryafcpxd
ABDqCzG5HlU3L/39L1fsXidTA2gCqg20YuRY5boIpVBtooidTqm5ok6kAbvL4b0r3wN/D3f5fgkp
adax+JxhN1LqbtBfNTrt5PGRuYlsCBlLi0ttDuz+8s7JPxV5Z19gkcPX7t96bnbwdAaLIbet96nQ
Qe7mdPIWkZoEhjhv+aMEmBVcHxiAa8NOjhQFwYfNfw1lUVqh0BRjpvE3jCcUetbmiW7tTHcOfZZA
6NM9L+vXQiuZkn3Vnf505IMA3Z0UHPcXXmjHKrtalEGHZot5lIWj2iQVypMdiXf41RqE8TGL0QRr
XemxPSw+U9lbQy0jDOnOSqePydh8W/QscflZgvLxfvOkHjuvpcQfz5RZWFAD6dQv1L06xXgQzeGS
p2c0A3KukcuXo+sOw7p0S0TBV+Tx824xSuveq65KOPnGMyXpDhzWGlshhUyLS3vX3xeKkNkt/P05
7tzWOLaQXQEuDq7DXa63fWu8QwsokyzohfvGK60l+6NCHVjogP470OiD+xdH0NuRAJh5MKNwwQ33
vglOFe66ErrnKeElLkloT7ZIMRUSsJEeCdcadOu/BbsrPmglTLViUrx7JcXfJBPoZk/cAdHl+T2D
2038mzBEP3pdtIg5F38RXVVBAjMJr+oZrdCYPitiILHnzRALBeBCF4SB2D3S8qx8PEzX0HLC6IP0
Ts6R4iNgSXeBEg/XpYVQoTutY8iUHO404mOGqmo/42bOAEhvFEWDZIcz48rQ/KlOidllcKcoNbTO
vma/fTf99+c9KeTvoXoSn8QvrYNvlq2vkV5iglrMZ3SgUgVH82sIykRyK4DxVDsKImUWHSffimCc
3qpZkeOa71eXxxwG7RrkS09otgQK+arXw3n0N5CPMPAliPdiLRbYVZKmNWez+EUhbfl/XUxREIia
nB4fKbQX3PNvRXbP/PF2zGC3LjUtkeeEqAfxkGRrZ/QQJAkIDeoMSroiqFopokcINoC/mxwbqhC+
HypXVKT8y6TGZTB4gA4YSMgreMldnI8TCIzdFkBIVfN5YanWVEqQWiKP9xttZq2+edrQPQBbE1eA
vBajhhXd93kus/g1i+H8VaNiaTXHM9OMgog6G+Ae+qScKvy5t4X8vEbVeFTM7eqjvAFbuZI3YAwF
qxkIhSrUFeD3WWgvqudB8H8Qmner2RYKT3HvDctSaORLgFq4viYB/ZyxrTrT4ABqJEY5awaX5IAv
eTdDwT4Fv/vJ8e0h+XbqwxmA112QQ7z6UwYP9ZhCqr5yOOWA4Im09LYQtfW/KueTyd1fZmTru4D3
g2gokaRiDtfVBL6CGw9eUzps4d/1S85wVGjhqLSrTovD6BfyTTid/HOcQNlT3tbTjMfugm/lNu/P
KtCkq0Fk5PaK9K8IuwiAu4uYQQl1Pnv3IqCatWN2lxuV52mO61AwcZdH3oNDtZmSfa+uDOPbVsPF
GEsnCQzYpV4+rILR28GHPzJnIY+2ADKwYbPPLgNLJX5HY2UfVTTxybYG6DGoU61+mgE0E8yeupvE
KmmjRDkZjo6uggjCklQTu+F/ltkgrCgS1R/fUL+2pRtssurgDBS6htGNeuFL+s8R6UtYLLv9ikHS
4OuUnQAG3EQFXJfDmCHqLRwIdTSrgaOjGkOOv1Ql5rXO125oTbiEpTkec6HY5LOcbeFgmUUDph0o
F5A+s1C8Q2s3nsNCV4aa/gY4hCQ+JqLKT7P08xl7rD6sxXJsrEVi990EwgFyyACQSWEWtVWQhXk7
Az6i91qBITTG9UX7piwVXScoEI43dPpeGEhk8/NFohMP4ZueA9uD/qMqETArGh3912JvOheol+Nc
U4AbJFg7VDsKCk97vlcf7+wlbG4TjX/3UUZzHHpL/w/TvT4XvZ8FnfdjB8VvzlX/xaC45ALQ4Q1i
uKak8VWQof7+lS+5ZME5Ko/fmqLQmDpQDZQyIk84QlSt4rJ78iNpZx0qEMNMK8CGw4vpytVlNUna
tP8paS3y+bFgpR03CECMklV3zPKs7ql5kwyf6u3X8riLSvocfhiswp2Kl5zvnc8C04o6aBEW/YxV
39em+Nm4pcDEop7V3np67ZHz9MSmfN/D95uwA2pgmq1ChWPYZb9XAE6w4tBkC2FNRP9tK8ewaySl
0QsUhNvhQwtZclvxuVhJzr2tMaG+xXSHEPHmoDDr7e279tm+GI6zSPAXfxXan7lHMCUwQSsMdiZ/
WzWwBxCSpHckxPdmA3YuHgKdLiQySk6RFMMcxRdwbKEXg1KG5zN9rVW59biA/x1pEljTRYaS2JX4
bUbAxwC7IejjUCJTeGof5yWqcJe8ycq7kioxTZyVeiuLRIfoNhiOxMRqghLf4Sv+EF6ULWDnGym4
aNY9fT1SXM5Hq191Kr2tqJTcw/BURoDU/fH+crwwZA7gsOqSLvkQg4l025nD/YSbnxK3/zId2+4g
1ICdZbl3clJ6/vvUP9AEylI5Umix/YcfHTLJjRzm0irA/DZDaWBSkS2QRvoMjUZMbVrwA8Oiuwqb
iTurDmWa5fJm2zcomIzpIlva2GLLIoTWhRMeC2+azTBO3Z+U+HocRgS9IIFZbLiCD9ZkN5L+y9EF
YcyIylU87dUsB5A0hXnXs14YvVj8E1hqBbUeF7gF6KlBHHEbQ5oK1NWem50XizC6ZF7aBDEulgpj
Te/ObHCMf9hwuZfLGmvPNyMCLZUqQessnGHY2iRg7rcSVoyUrWP3drY4B+22ZC6oihuzmWa72NoO
yfzdGa3IHawfC0/9TaBaE1ghKPzv/DGA4beoUSuc0rpPFsI6gR8pxFSRmv5t08vNRc2wEuwbRd4x
8TgOqr93VCLI2Sd9OJFyHMDQwneJ6Ba5jlTabXjwpWWdYRtRScGiJeMQbN8y4/h4XqzOZ6jktH3P
VXG/2ZlnJrOQXmVI4p/5zDuD1Oyzy81/XjEAtIlnXm80I7LAOIc/lRC+gJr5f157URDX5xCRnPUT
KTEw9HVz19Nr4g35XOGVPrgaVIu8/bRL2tpUCvXsNfMyJ8bOaPk1Kggy8FpDzPMhcbd+HQuJIO2W
Ky8ap5GdGPSPS4c+RXVHfGXFt/GemwpS7fhNGAXJmCGFI235SbHD3nMoXIN3F8L1prKYte/vI+DE
mVzxFvoL2kaB86AG9pTalPw0rnyI6LaTRpZvSYG4oDbyX1Qoj31O4BbBVGd+3A/n7QNx+p1n+DpA
uBm+S5EYshohm5pFQXb/s/sTEP/DmzstwliHZFPGe6gDGDF9/waDFyzgE310d620am8MGV9Ay0oD
Gybt9nGuDgWiTvmk9divQ2aTl6Sz+VC3E6ByjEiq50v4Wk5dMcjpwvwZ9sFHVNEj7rZ4vDdWagEf
E4zMRZwqhUw0RoPudgUeBZKkhJzk/fJ2grv2zo3vdYEVwDhYFk2sDED/6ZJDqXDlUPm8n2pYKbry
9NcJ8FmSi3s5A6w9P8kq7LrNVvVKDudbi2wAq+JSLpW9XEQNLoi3aKVv9AipVlJ7gfNbn9sUtoJ3
cEHGY7NBSheOnsjF3v1FKA+z7rhD3yT5xjAGcctRIRSKMNjlYo3ggDGuOB6EpzlJo28Ic14WBLDX
1ZIDkqSs0rBmbN/mSS3jDozzND32MpdJcTgSjzCGtCfeTe+arKSMqMoC4aoQY0ftkPVxTzaSbnja
FnSxGa+AIbn/+xFPs9PETgYuoo/rbf62SSVeekDQLX/wuz/vixP8Suz1b/hwXve1kjP5PU+qPZAo
/iUoOa3tqxRbaifGNzIl70RGMIhUuXvgSgbkfLiJb4OEsboQHEVabWF1knCIwfVnN10Wg1iHfYBI
UDVPPEbURID1iyd8uNJ7fv1izYZNjr6wz2gbp6B3tkSl0zdSRTgfoZAx4tYmPJLjHZr26oIzr8L2
3iPhcBXRUH4jc5dYLLLU3YHDzZcxM6B/AsPjed5x6pDOQJwTS2xS3hhQMvKTwcyGunGiUp8sevOf
ZZF/jS9LoDkj4BRVHhI6xayLtwd1M13cG+dKTdrqPu3x8QnaQRYz1LCq1eW1kMVEiJ5+AjE3fbuH
HsMmSd3SrOzXpYm7M8WsoTuSQ+4RwXKcNpsTYlueJjcbqVAZ0DWOJ4K7SrwVb7AapQ+Xlt+Pgn/p
nujuiL4w0MpIvpwMzcePSIGVul043ejy8w56Y9B019/VCxGBCYr26o8bn066DZV7MV8t3xntBq1u
JrpgHO16g6QfHQcvBxxOHBPshIhdEtd31sFm6+brXADvoxvEpW0oZrIwbkPVxwOGYVrW3s9vjdrL
oReL9yQ6/6GTeNDmKteIWTSaVRqS1Y3kK9yKhr3/yYeBbUE8Kf3ybORucLFHFzWdyBhDuKT8KVQ7
gdMBPh4RvHjOJlaZUmNVQkuEFv1wi1oRS+sAfwqNAcv3mAEoMo6uvUqchvYlVPpzUEM9KqNvu2MS
7ZhkZsUyZYocBLu8djKXoqY5V9g1CZVXTk/psXYV72N4q70+9VIhp7StbKv0Adahj3Z5NwWUJvrs
hLqN/zn8YqqW2d/pubFTO9YL2ci/r8l6kDyZW0NcSHj8tc0H3b0L8jQpP/jFYInrPK4dGXp2HQF+
hrI+jSv8LJUuHGUuDMhi7orl41PhViu9/gGmGXcn5jaNo19JjE8rUkh/VMbJt8R+ln6lPDIMiW17
BAZFZpx9S23TruqnDTtoBxb4ZoOaCNAgu65EjZHtXS9pRqCE5kbyGZBxsvPAKBDpCZK59xd3PGuz
crYbQzKt4Ahk5tyuQ3qZvaVePrCgudwof2uH7f3vckT9aSvIksCmn1jukMl+wlpEr5cvkZV7gFm8
NBAJ/YvfOFgaYXMzs05/Nn8fHZwZ/cQRxJZSEfMYtuaRUDRGE6SXp/f9POGAqcimXkzdjOn7F1YR
xDUPecDwDNy0oQoVukyUtrTs4txJmb5/n3ddtknoCBo5JbJAKD7QqmQgxSwk7eSxRSItwenoAC6V
lYcei1JPvaWxbz8ktpE9HPXW9U95QfcyIUpMKOCh7xEKJjn771ziBn/hZIt/p2UXSo2uRTggowDY
wDtLAE2xdsXzwevuJD6toIdEQk2BBX2V6e5ERz8sb7tL7c27p8aLnEKvCqNgcVEKVLueipKlHGno
G5T3TnWJ05eHgBdtA0V1euA1xJt0R76GZOvagTNP9I/YetqWt8ZYqwF9CeA2boXWb4L0Fvx5vlUG
5ZRYLgKsWYCraaGKS0+GVph0tBVBQUBJPtcojyjL38b/LWketXk1w4W8S53jz/USFxkZbMg4me/W
I/b/ojGSSMnxBdmY8ANFQjDlFP7ClJc7WaJmSURce4B07zjbA5zqxNmNzmHE7kIh0XwRi0c4P9Xe
oaFOu2cBxszub2T0BvXt1RWFqhLIy/ix+241JYLowaQMq2JCY6wzx13+PTgJOlcSAh+x2ktAfnGX
E+VYj7XvkzCxXJqb1WLBbaDdUWXnOCUAZxgHpVANFmOwXJwDcYeQvIzzVLqcyK8LqNpZ/IGuRLHh
4Exw/3+NqJeL6UaV632/YxCFdERi5aWVmc1F7+FUVLiXvhDN6zJxM4Tmk1+l7y7zexCI1bA/Ktf1
a8WGcjmiAo6Xeojf/bPkT7+5zjF7rAmmOTHCXf8G64BDiWQbihWrw63e6J+4nL38vRs7PEtMx4PR
gEXPhPVxcUSqal14mByz8pOaJC70bgYFNyYKScwilCAV4GqFf+ngZyYSJIlsZVvE0eAzY6qwd5ZL
4NhwGWkKB1v8AC7LdaEW57A/JpYFg7TUJRtSkShqxtnKT+nQM3FjTOxvlyTYxsPVIxk/jOw7dzgq
HZ30eCY71/1rkggS/oc5Q/GRnH3g+qAA51GFaVsCROqEC5AZSQaq1y4s+7yYAQiWsg1jP9uMUPsk
DmgCuvi7nDxS4vdZzPXss2PebdnDIrNlNAyEhK6+s0g0uCBhm+rNZE4EjVLIdKa7xZWbbgv3Euve
9qolDpUuXFrEW7eWutLWp4FPVL12tnupcGw1kySu9jywrtr4JMDNdSRtdC2oB+oGgvfDal8qNCr8
2b9hwwH9VxlRDUOWM0K1V3jnsqXz/4lh+xOqqBPyk+d0AZuVrCvJlOTUqcwDRx5Z458DJiCQYHUc
a4fjyvwK/c/GH+uq9WVXQASULiBbrsoLcxzDKaDEudeQb5yxGNFyZuf9wwHtARXq/sbdOUY0MUNY
lnzsT6ry8tJhThA9QaYK8G2i2pwjEWms7gGfceMzpIxpEiRCGL7v6tZAGHDfgav0jucoolhI7NDv
o0UGtliRCkwZALZh/QlkrgPdstcEkC/FUpD8Vl519tPf9YssGaQg5inL31q9RWlg2ofqutPKH8VC
H0mk0WAO+6P2EaZOczWZezKJ07DTgfWhhbLa1vCvvNq4BJ8byyqj1ohEch6RYKKTTMkldK++lGg1
xfwCfSWtUazFfnQOGggG4CaCYAeHM/pu1+hSedhOkIQCMEeiQIhnDnTskoWzakdQWYaz9zItp8sM
H8a2nW1It2U2i7ihMggEoRW5Uo6PJHGYei20D2sbPE4HNzswEvXVVANI/3fgOJw1rX6G/dI37YnM
dlBc8A9DsAOCQJngYzi6UGNh6BUoqnO9lU7Ugj2TnNSNSMEiyku3C1eDpyndYWuJ88zA8QRCcUYy
SOWLVMjSMK2L+GFr/xzUR6Qh74m6HZukImQuQ/HQBu2oAND6ggR0vb7xQRzhhm659iIEdoxRCapW
VyMxbcJ7f4AqH0PHZIsthw+N5rEgd+aGxx4kkR5xSOOK7NPbmbuUXnU4kBTLBTqXhMPUlkxZ5IAc
0EWGB3jmmqQllll8jC1/es8xAUnpo4DguqYEzptHEB2FUp4qSuF5q335/4ww+S1N0J/rAzhmCuZ7
GqJzUxqv4vURjfFSKTxB3SU1NTQbrgV21EkXGmMzHeRYo8R3QV6R82lIBwrp/sAvksljqhXZbDZc
DFI+2qxSEBKjZFXhpIXzLJlDfY0c65teaHWBYrNMCjjXls1hnjOTA+qJXuwwxMLHPoqtqEFi4xGx
+M/Zl8uonE5r7GmEcvr354gFL0iZfPrPOA1nFi2zLrlLeUNrvnS2QrjDIrulSJS5DhYIs2JDWblS
IUWvaJS5III1jdVDiZzkMDg+h071a8B3fdf2+DOGA/FW7gb0Jn7rflez7xMPV7mXTUFFm0xaScIn
kWiEnStQXGwHtPzid+MFtB8bP8b0XYNESGcO2g0EFfg6143DfHmuPyw1SsqSiunsuP+3k+5Awujf
xE+O1yTRlXEDnhXzbWmQ0vU6yCOWx28JKfYYAJX5Vnoh1Oc+P+/cHFqxr3a4K2yPGQswjr/jC3tA
QBOdtzw/fym/bUkjKPBPD44zFhhN5owXr8Ooh9zcAzQ/2fwUlBeRW8yg8xf7HJ9YlQe0whqHl7h7
SPtRJbN4uwmWM+VRR7WAeHaHfaK1J5AS2DQJfboY+SKNNdaHosNyiTFS6MRDbifO56QPhI0G6pZn
+6tjE/CcuVKiOupz0YFfV4Ou6bKUZY0KrpXJQONPCYJeta5TJwVELC4hnCR671lTZKLgXKbRfCaj
BdZeDzpR1BzXtaKRKhaqx9rs+vk4F7RR6sowox7fkQPLiwlA0mVQb53Uf8QH+ZNRln43rd9X1ETl
88kZSLCWWIceN9rK4g0tr0Au3wRy7/22623gZMHyXF/92eRzuPPS3pEopJNbdBeujw5udXbjhZ8/
QqD+MHFf/ATyiDR2mgrFuytl7WvTjioJWz8o3ftIBI/SV/5oe1SByhmE/61J1QOs9ZnZZmH9G44N
ubAMZySnxxFL16cqJ4tt4qUzqC8/U4+xX5UnsCNODZGNpb2S9ePrHv11U6PSgjH9QYe5E+CmS2TL
ADRmnwMxqzIZdwoA6rg2cQoe59yQb2hdWrSws2ihrdBveIaB1H8IQVL8nUV+UGy0f1SDvCE8gAav
FNgRuNf/MpQ65NbIGUT1JleRAjpAGCYOFcu+z4eh3TOQl6A7jkF29sGTi4WJn5loB75Id77tYrqv
Omus8gsR02s7NP/HS3Byn4ZucguOK7nBToJWzcUFKt2t+w5hqaTy6WeRFAdEk6Mcz8DNn/IGpk1V
5vMSQFuiyFAxFneAEKbrFd/vMIrWebxqNx3sB32dJ8g9Y8zpwyiPCK7/mrwJr5HCqdZlxflI6rU/
M8dhtTSPvYxpekdJe2WhzHlbbR4Lhp+XqU0eI8kn1ePRMqc70Ozc/g1lr7uvBEMD3zYEBsvk0C87
63HqerJziHUSMkNOxPGchQHxgmbF2xsRJ6TvlaYZLt0C7L7JKhL+acIuJSFaHw14B3+r4kYg+q0N
952zzH/1jVUIoqJ1wKOt5Z3aTGmdn19UyZwd+CzxFT14iHHkmyj28AGknioSgEbzeHhiLali4ZbF
ce/ozdQRJA2AHilgb0VG21Z4+vhqPFS5KQI3gWpL3iSDOf4vokx+Ean746xHJB1gQfHdp/ZKCOwH
0Zluvxa/EH3+YlJe7IKG49pgsiylMxWB9BTpR/LFDBMHLy0fwGV8Fhp/KSeVVKEBALxmNiRYSzl9
4yF8WGMeLshANYimQ/Lk9HYjuqZDQP7gH8EiVGrLZMnKKIstmVKxxAoBvhj1PE3zPQncGXGZur6o
hoFf4C/AHbNx/T6rv8igCvLyMUegzpzQExDRrKj/BJ9L1hzhCTcFx0DoXLktT8TT7tT6+S2ITCpb
zdMBxLjrCkxZQRZYFF3GZDUHI3KhQzzcDPX7euD8KCLOQlHZH1FLcYFdO2FxyB+6lLhPVLBNd0Dp
HS1A
`protect end_protected

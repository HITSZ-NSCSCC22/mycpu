`include "core_config.sv"
`include "core_types.sv"

module register_rename
    import core_types::*;
    import core_config::*;
(
    input logic clk,
    input logic rst,

    input logic recover,
    
);
endmodule

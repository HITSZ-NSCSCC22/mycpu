`include "defines.v"
module tlb #(
    parameter TLBNum = 32;
)(
    input wire clk,
    input wire rst,
    
    input wire[] asid,
    
    input wire inst_en,
    input wire data_en,

    input wire inst_match,
    input wire inst_vaddr,
    input 
);


endmodule
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gZu1SY8CK/JrHDtzcU8pxbpsZaBRTduCD4cOOcs33DtfPh13Z8GDRXffarzKRFrY7wdR05orYRHo
gxz7VEq4Mw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oXCESE18H+hgpfL49akiQIfn9nwcZcnlEC2WeOVnRZujDStuwEFNLW8q440rC849j9QGBfbyDMyf
PucktieB2E6u+IN0LgoXJ1hviWXi2aMTjQwJbzKI6Y8s4VPtyG84zwZUSgw3MiEAn1ND9wZNlsAa
5SpZn1m+6brrdKttyoQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lDDXJQQo9YiwNTEImWd9UF1if3cpWTjubZDL55FHgE0eIkI2wz5HPpNQ/YoDvayQRlzGQowduUVc
KbxReNKJF8xDlOw+rmB3+fosfILAltXM4Je4S1PRa97Ycdpm1ae4gFTSJbVzIvOabZ+T9YUOchsK
YatrXkJaOo7JRI+ZJhMDzSFFPx0NDqnG2wAjtaGWMYcQYOlDYaIphgVdOOas8ymx7ZlMIFw6ihK0
qSqsc40DYmLWa2ScMmR+tvbZt6Gw6zuQvS5FDfYFZdd9AkB93755fbElWNCmplvCGNKSiUof4kyn
uTTn2MaxY7145LPzLnJ5nV3L05FgB6ly1RgivA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kLGuGwC6VC/CenJt4x3XjzbXlZm2Tsr/XfOh96IXIeIUpnZtyz88fWkiuR5lEWmQd9O49pZO+ZSM
Y7Uzfd2FzAPCBgSgpmfTiogzFeLhjL9DCHKWixiWCrV/3LCFC/PykfWFtKkHgVRkgIaCkKp+OV2Y
O2g7vJgLNmUUz0Ud8DRky5S9ZdNddTvjp1gVtFMc4FdVHq4XK2jJSUhHCt/0wEGsjwHkbKR/NYzB
9VYiGjNNDyn9G7h/+9BKp9X6NJ4o6cpBDvtYOHMMN8vxhdpeXpDQbQ2ZCZ2FJ6///W4pqVA8cbUL
jtHfXmYh7TSwmqWAQ/8SfUezLv0dKnMAu4jWPg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ABRUWHDQKJmsPu51jP6AsLxdDI6FEgj8GdIFzkrmZFBX01jO38w52iWwWJvmAiFPGX3/jMgesCaZ
36fkKtn/zf8h6LbOffuV/7ay84ETINplaMD9iuILjsAZAvgnxUd6QYQDiYmj/Nne3qEwfx9Jxz9K
YJsJn+iFfHbwST7oExnh0r/a21x2xnF7st8mcek464JElNN32lshx7h1eGcnqVdjpU/igI4R+yPl
7Ayw7qiaKWKaGccaRrlJszfFVOpAyv6WS9A2Iu+Doayv65qg549fhSoT0HD0b+OjkzyFZ4xC8aFa
OFSvcZzBn4JhJYY8oH08Y49gKbijxuWkRblkVg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kWyfC/S+TFffzZhIxHq6+qXTXdobS7d4GBAW9RnlizcaO7HAxuHulghCua6DtlcbGoP1So9G/DLr
kzw6K/IhnQMpeB8wAhs2dqFfbbGJvNznLIqFfNyKsC7O78jPw2nZa90SvjPoJtiR/LjYfmjnGqyg
xGh3UXuBqTwEB4Lxu30=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
muRoSs+bdtmFFGZd10wl0c9URf+3ol7CQXPpbBl52a1hm+uvHQVoN3MZZdHKGfqX1JBLdHsRLQCi
hVB8QQwGUFg7nSuk/rGByi0cDLUcOLk8tIamKjJemsA09GKAXGHaPH0TuR7nxAnQrKS58vEqPL6+
ibLavPNjrIQ3UEH0jji3MXKRYSTb3BU67W2MSVVFTgpdOGL0IF1ACnSJNEE9FJc5VsyajB5sUuQN
vl+aQ8OcaETzGbQQeBpQuJdrgi7lnuLyRc47x6zrAIKoishoCGjIUvVPMQZ4JdCZCLFBphWIA84E
YwKTl02iUpY6G/Imx2PcSwrulzGAZRyyT4SliQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 566304)
`protect data_block
7VP8gCnvWMaXM4YnOaex8GFJZwW1FD+LMYO9z//oKRCT+ctB8KPjfwxpWwQAe/N5nIpX4khcbMKo
wRaYAPNPZiGUSqWIjvSfQ1e1y5skfGCyuwA4PnbBnT3pbx7SW4BYNnezlINjEEMBj5KY0KhcEz5a
qtWeAm61YTOUNdi8OLCnzQplyeXvEXF6xBuKxbE447L6Eu1Lx8eeZ0iBchHIkd9NEP0MiiwUeMDX
y2Yj0UEBeoJ1Ea6Lx5PZMmDS4JtZgpFjwDpEqeYevCzAh5xqBqU/oLzcj34XoPKQSfKwqChkrv7T
Usfv59YCsb4nD0SmOHqiRwzDqaDvvHsonuYXXXS4TVTvRrvlgydRd0pymWDHfVY4hVXYpUKJZ/Vz
VgUNecf4wel/BYvYjhqJicVwzdTwwkJy9Afa7IhRzVgX8RtmHjGvSGvBDQS5hhrxhAvF/PUrBfpR
2CXqAdu825Hc7SRqAef767n8FBa3sZzMZcqk2rlwIykpcpPiZSEs+XF+I7vRbPyI7um68S5rtyO2
lpX+YZGx9YwXLXP6ikw2D0Asu7eiyMeTvk6717p2p8QNjB7arGz+1fNLWUzrnaPtX+JQxuXi4Pc7
P5/cLgvtXBG/E4AK4xvKXnM0On+EbYeS+A7Sygl0hgUcr8OdwHumD4Dfhkq6lFfjlz8Xl+AIIIJH
OBMgN/t5lndftSe1JP/OzOKcfdRexrjUUDweA78dl+C+yjY/XtRusPVoPkOtzniCmELtklpGsL9o
QlL0yPn5S4gMqBHpqZnp2HMQdQ7rAk5jU0hBMB2mQWCaF6zh9lQnM/eCHfmyVv2gzmFsUWTiPyAM
gsZQmQIop8IuFOWupJ+W8WOmimHcfr4oVX7pa+hT9WK63kJwmvHzHqXkSED2xHrMREzJtirNYERi
+cZHSQsNskJOMVqDx9j6TcyKxG/9pNf5Ai5K1EkvHwWl7e4QFFffiZHrbN3Qr33wJtTC/+LNi3rF
qDVz4QGQegmUvHktpjwzXdt7xRmwVBBN/J0FID+vWo2QAokF9KckmeIH7PXx5gYtP1Y00yjNrT7G
4beSTvBFCdYIZE9GGubVWg9rWmoXWfrkujAoJATzbsh+kqBD/AjEXe0xI43U06anKRUKtroFUPLT
DQxAFL1nRbk1Tqxy08vxDbItZci4rwjq2SsPOpCyV/LpOfOEub2kzSTgLp2WowbuGa/JXa6h594A
yi3lN3+DBqeQlH7yFNo+Bt9NHxCXnt4BDj1v9Ns1ljoSdRjm7Nyz/UMwdlvTss6GOrTe3EsFCmyk
MVrr5AxWg0IIvLJAnMkqRsugoYkjQDwAcym7ndB9I0WdMKMM3kEPHvlDRdTU10VLlH8IIFIyllMl
D6fdq3jWrU6JrRGoM5F9m2l126yij4jB/2SZclzK858imMN0tT5r8qjnsQQTlpu2kn278ET6/Gtv
jmFHterZ0r/2yZNcNhOweG3nItH5ia5Bqg6A3XJyNpxgZX2CMindsA964+Nj/EQaGl2COYDnN7KI
jVp+wSMmPcAsuR+SI38ORAFzDcDTswj4gnaGSRtroCyTmTvMuf3ILIIJgXtdoIpxdeFt33cDqaxK
MhOu+JipcOz/4Q1NfHzssDWoL2VXp54PBnVqXPfQWNQSrC60ksAHYaeS63kbMIjFZoPHelqLv6lH
/NJgpGYsMUVVwEE2h72j/RGp0KahD1Pk6bUWFWgD/ffd+l28on3z8ESvkKqV99mBxJclGFiD+TZj
FNQX+J+NLpKXCYoDtiAhPke8Xh40XayfmRnLEHYnreI2vFT813fsftvGVv33o7EUbFbmSM40jhRo
WgMDEXFfqCzJKK+A6uX4yQbNFzYupsAAO2rr3w8xkzotfWJyb/CMOrpLMEQM0pFMIdMibg8wssKr
G5qi+O86ljFQGKH2kqMTPDnKk7q9TWhGDmjqmm7LvIbUuh4yMP0+csJ/1AECgsiufuqLlpLQittn
euWFD6Knrn863NyE1EKX0j1BXhlnQPgape+rEFnyr0zUG+/Dp2AVpA99umsVjap3ZsO0x9KIyotL
4OUfNDEL4ReU1/mEeJy7JRBpBM0xoenSzdzu9L0Hx3RfBPDBeU6K5x6sKf0GHRQtb++JMQfH8dX1
bsaXwFroXQMJaZ8/prTFw1q3aMv8iLUYRfim8kUfyRgcywvhbgO+CLrEUgp1LOvZ0qVl6Kqf7Jqu
2ZxbF4OmVfVQ9xLVCZLeunrzEdYJB1XmMZ8teuRBc0UON6BCiXbP4HToOVdsp5r7g/AsvWV9+NOk
DcH0nL5e8EdgTYrazWCGPpSG4V+UYD87Cuctq4ErMItLdsv26VtekLuxfB3XPuATQMnMrk6Eb7Qv
bsVSBndlQeZBgLRzMM5bNiB2xKoU/G/d3hAQeO7HHzb/VLj76jkZQLNHVr9hxCO/UfcnM7wjvd5q
ZlGBsqznrEp3kthudRYAOd4xNqwHjKsvkWJGgqRoRSC8VrEFL0g0ytDN9i0yz35ovLQ7FbSbJy/x
74DHVreyXr07LKpEnkHAD8NeiT0DZJNpQruhpNF6Ot3YYsMRi2KkblwzRS7NbzuUzy3MhzFSykLe
hF5SQEnjzpWKEeK4EPeIje9dwrBKXpQ8OxHt3/mRPukAjAY9trdDnKLTa24pEkH5tQVyboazxoEh
KfH8sA+cD6ZCBKAKsw9h3j+Z3MRoNvPDid3ZFLpyd8k2cq4M0dMh6uK8HGLTjeH75yQ4U8eC9vr8
/PUB8IC9wIQJx3QQ9m8rv9KS3Day63EMMGLOkIf5124MbYvK1aD1iheh81CaGLdgTICJzfNxxetA
UeNP/NjeB949yjcj8wb/SrTnHmyLSx81sPhsrkLBFk1WPRwUjUZiFZVeQBsSUn5KPFhhddygmhrN
ZdzeCDRScFybLHuhJX4qsNTAIjlFQpR7+BM4zyO2/bDS8OrcZ4RfzFBRyNsxl5KXmqkYHbAcnGMf
9jGMl8KpyNs/KXtIIOImMVQ0nFWtT9ZwZ7fT9QFhS35FYy84CMYrmPC2lM/VyHtJRWz9UB+XMqKX
SwiKX4xtsoW7xZt8GrXRrKl8EFpzjAJHmcytEhMo1bJMhbIWwUmHk+RfM71IHlmxNvlF5RBiGSPZ
rzLbNBt51Inm0dL7Eou3slbnl29aSEdA0UxSiY8rsnvptXgwfNE3n+4GjRGfgvsHjMsxQ2ErksXx
YtaqFO3F6iZIn+tsIlk98Lmwil9ggLyDlWxJU1C3fGBEz+eTw3dAW3kJvwROFguf9XMB14qVhaHD
AZhimkY6cZVt+cphekUbBPXgQNRPtumayQvnUSqDzUG2QmvkaQbQOOXWRA35zWH84t5/xnMZJX3y
xoKKUSib1GYpEodsGWnfME1BQQFVJZ9KrXuahB1Syw1wO6N+VRgh6l9gD/4WVck9T3XELwGGziAf
iQtstTexGgq5FRNOJtg8kw6y3wnyDssrWTzp/+5w5vfLy4ap33pfS2p52czj67fOPKqgpsqeyY3P
tjV3nJ/B8rILqrWphpUMYJ+PqFNq4iqDuBnHXIXiGiSJlpxELBuKlJoprg2x7NQBJLSXT4H1PgyN
9C7xrEIoC+0f75aCKr1AoPci+etyPG1MF6+QjvDrgF8QPOrb0LrjMfVFCIWRnE5mG5PnR7B9QRnC
AX1tum2Cl+yM9PqwNDGvbrcNqWHtHpTq9xpwRlSdAcpy5CO5rsCVB/JS0DWXfMf3wZKlB7lVyh3w
nLHRAjt1deo3eDENGe8jiPdsmNqHDf1+lXRYrVffFXHbQo0KIwzl6AnRIAjR5xnsDfSkbqZ5qIW0
/33P7wOgntwmrSOfKqMWuKaeFtXOEDPFDnT1vy+KcSrXDmL02qu/R9zgmobSv3cpe2PqMFoCFAa7
On+A96I+aEBtj3tVvRr83bQCA+v7aIyYwe5hzqUmE1dvYobK34pAJ9bKuidEnTAx9jHAmOI0/LQD
0uhG3b8gte79kc0hSghhOFsHORldZgZRfD5yMBoZ6Jw291pr335vteS9XtEWmZAj8H9s88Q/u8L3
IHjIQF92mV6QfEmN1mzj6NDwP816dmI/WEcU/F0n1SWBKYecocN8ns9G33TTn3p4vIpdn+Qwhq0P
ajMKLQrL/DonW2PLzYhVy5jPnwNEGe2QPYY4ysgAq9DjUhyH7vO+UrtX8KHdeOKK/qtrAAtqVC/a
ef/Ipu5eruam+yXA/cezYX0Ahc5vmMqhbIx3empMm+WR5sOapPUHTUm6LJQrspnonOWkUjQHEffZ
AM85mOSSyeRslrSANDlNXkoCUQ5o4h86ThNF8As2IKlTAvI/15sbjttyjPGZpil4+ckbbXRSjKwI
XzFbf5xWQ90IP2MEIZtCqX10/C8bFFRMvKvShmS5ouTr3f9lcsrrfHMLFDSkwJe4/dRIVhCTlJ/5
dCSEQNKqz+TYaVsn+7BI4cJClx5WEe4uBNGfftPcr+Oykw7DAI9hbLTSyKmIYIhF8Wzvks3G3RNP
8icJ40GsfIdoc7MengMYyF60t8qyulMJO2kZZMBOUnhxc6/cicFH+rjMmuuzote8hudWN25tKg08
E7SPmwqgzcsARPLwdG5/xU3XghyaVWHDgVSun3dTFgUZ3vbh7IkXfuy/gMFAY853IhEaxOR+DasF
uXb4LtfXIVZD9FhEaamvawfh2+Vztk6YSoSh4v7Ekkm0SydPUWF+l5/HqtNdEJQyuDGmV7iOGBwC
+BSMXQRvi3z9eywGtj2J4Nk0ZAh4i/FQD6yeAlyXHGJE9DvV65M3g7kvvuhGVqCyG1Y3GkOKzhS1
8HWpM0F5meLIIep54J0UvwzFN590zDDydOkREO+Rdv7oxNU7pZYWfr0deI5k54/gOm/Tf2LEFUjV
7pAdLUb8/rqFfBYVOFWVYQjcejb5D4V4Iwlet8cuOR50UKEDJMeSQdFTy9/vYFS6QPt06L1aBcTs
+dq5nbCqZYMn6rHSLmsQAyfvWt35h9oBCotIkzaHwYVcZcY2ePp4TLZNAGuWdN96p+yVe2MJinWx
EhBsG/GABP55Jmo4qE0Fg6VxOHG6yeFw+9GPyQVczuZKX5fg71wG4PbModvwStaqK8uvyExsmWlZ
DeIeMYLNM/WXVvv+lQ3eV/cCufck8weDE+97npJm/X+3Sx6jNycFBdsGMmnuN3TkxZFoTKi8DeR4
tbyTnEBOC2QLOOIvx2+7JywnB/UGYuFi1sEi5JJfotbjocjpSVh6P/+1LYdA8LgW4kqNrY36BZhY
7bh7opjwKiV77AcRuOGyoAeOa9ge5xYlTfeNsqyCbaebqEmBl+gRPIbIizbNvHly0cGYcdVnsXp4
SQ7y9Xr+xLPRfdSJynXO/HasP0ry9g2lL8YJUOh3w1F5XrCaIX4wXzrh7TyEEXz+Kr5nFwCWkquS
dv4kpNpWdp7+ClbpYBiyC7FHxJD1h18cFFS8bp1SMuWweP777JzrE99zT1IfTNCqSb2FmsmRCKCL
kFfjy5JfSvre7HU78H401MCk9XsoXbC/cOWLOJxlVSzQPIFVuHxeEewKTRfJBXB93WrQmU2WnNAW
JhAejHLNjvesZjOtc9e7jr2XDSVPJw4LAD/StCD/hHT8SUGjSvge7e2d6a8T6s3bY/ycuNWe0xDk
WtLJAttCjnP9oQu4dczlJlsOJ491QPGuwYIsXF/kcqk7QwmEi0mg+7nE+krAKSEHmJREO5RR92Dv
uBJF/jo/erzmEkYyYWaBp3DnCGb//zATbyEWDiZn7x9iGis2v5C/kYDiGy65yFWrhnKT6rIfWs/p
xrESc8Xn+FdD+nBneLNAyDKW0D27JWf42mZyBWjMRxsn8trJoUfwC9qwLhfB1/wAjAHSxx2jVypH
A9wPr3aTyXeSVzgREdAdfQnKvIYpieIaR874nLq/NPxTunmUCIP2e+yUY2YZ+p4NC8v+ubdLGGCc
m9509aYruLDvzNNZd8ggGELN7v9DVkydcAO4nVuSPoeU1Wg+Ofn4gAaaq1RoeFW5uOVctgb1yzlo
CLC6iIBa+EjYrPW7mBG/4mBqNcbcdpbKHp1VFuredzxUT0BNGmJ+pFCwL7a/rzg6Q2PuqCGVb2BN
a0AZw7H692vJmeZTRMn/WaONm+uUJrrs8u5Pb32gMPB14l7Iz9ztl6nrDGKFZRDpNsYsUXYey2rf
vc/EPpI6ttDgbt93ShZKOldiirB4JvIbESjedOhfqZXG3pEapAADmYFAjnUHdCC1jjC91p/W8Dc+
EdOqJGCAR30Tm4XUy7ExO7F2DzxiPlqDDUSfxOd4CYioTNhy4IIIf2DagA8fexjxvR5LkiuvqbH6
cvBsAacqhDD82kUPFYgwK627YuLZcMbNk5Wq3m50L424GEnWkQVN7W60LPpYb0yH7z7R2ne0FHTk
95RsyYBKAoUCHp9hDc5Q87x8Ri7makW8W8qCy7huiNxDOyQ7h1BYPkhCm/T2vKvrNWra0g7PIhTC
norTlEvkrO9p0ycqL8V1OAzJ0NqEJyAuB2XMKaGpvoqKCz2VtTy1jCnp54MMP/4gKgejJlx4QqJT
8RL31HZRWKQ8Kgm5uNEqFrZTlPe+nu4Urki9zvUCcvwNGjBt+kZTh9k7yVLEsU9qiq1NSJV8pRQQ
qZ1cNXHNr0WsFWoiQJlOEoK+jV6wzLjzy2oLyNxFQqLvJTY3u2hPEqR4jvhOP5dc9Kejly/qbW8N
kyxsnub3wjPTHyGd45kmK7MnZgdgWtl+kMQiEKKB3QntI8b3y6xMHVccMZLbnCZs0nt5HfD2Kgt8
xfjQRTiNuaob2a2+UMXDmmhgcRVRl5htJCP52W/uJ1U0VdlXD5cQiaA18iLD1WNuvJ7dwlP/84E8
jmGI6Nma/+Ha78vtqyCSUlDYOefl9bEpcfqAhGf8PW5+zmmueINUq7GxdrOKVbH726YmjwNeofJM
KRKjVGTd/rHlZHLSQ/OqGTxww0AG/EkMbPZGpuxVAHZPU4t0w6seSDElF4w0yXcvSm2FPEnUQYwy
izpAYoDM1jNUCswtCpuLJk5UNO47hxtXqh3CWZRC1mmqyan7UyZMFptLEhQ/VrSyY5sl9WyaPxPq
1Ww8liXAJjwHznkQVv6Sj3eg6MmZsJf8h8CTsNx5/9SZwM5MjvsP1+ZMg+rzAH1rjmJdDCQfWZrv
K2DyEaN7p4lsN+AIhYI67tTQPtaiyUH6mSLnoKXRP2p9AurGg04J2MunZyMbMDFeMgmyRWYn5q3F
TKZJLKPhqyjf/yI2sCkY935QLlyB7Gn1y5TzW6+Uh18v7i24qvJPvWbei9L/lCCFWHvg6aSPRJmt
ar+EWoIXbh4GWlYh35sh0O86trFV5mC3P0nNbPGyRYsKO5GX07DMn5rYhluk3q5mbGtfFKLzVZqj
xLBHWyDQu7ynM5FfrsDGaKAFt4cryRnCt2QPhjnSi4NJbUTx52S9KzCnV+MPVjwj9nXCxcjWTDRQ
k+mtGCgd8ufj2BUC4vjYnzTCVkvb1L1ysNarF/48sMij/8mwKAOXG1pKPP7gqQ9qUVrf/SuEwCqd
zbzlhoKM2RB1bMtgAfYmWVPR+VCXtySvMZzmQyfioonADtaH0CPhJzZohtqdEylBLsvW4TNLTQ2S
g17qzzWwuUfhKe6YjgN1Ck4C5Gj0NBoNVQK8kzXtWhKqxURARwqrg0JHPqEcEhVFRYuOU1zTr8Yo
32OmztEbgRqnPHo2Tiqw/SeYQofwPdPe6SAv1o6SuFUwOTulGg4niunAhEYOFD4iufdcfQ7wvAnq
hBjkjH0HLc0MMa4K3xZ6YId/hw8+JcXJ3IU4C3ppy2/q/MnOTlMBMUJ2esgWSFyjqhKeNzF5HN7R
pl7+Af9JTllHZ/TDgrFGUOXcFI+XH0/9ibF3V2loSvvF4u6mvKyjcYtDt9cuqCIHkrFEXKrTM6NT
5S4NgJ5EOwwTBUuRYi1EiKKEafih8IAcDDQMGkTavqBT/O69WeyFyxpXrYz0hJHg50GHpk5V5Stt
wwVkCg7FtvoKbJc8HS9RKYveojETxscr7gefq3f13C3/j7ye7MLmVl4H5yhiHyEOsqrtMgX6w1AJ
TVti18kvFRa94bExzOXsSa7CqIKobfyVrW9QCsxFDHH1e61NxuJ0egLE7VphQMcsjzj20qfbcJrQ
LKCtPBX0pmMsk3T0yTlWZapwJOqyKQ56qf3pUqls5b1OEQVn6tM8W9xL009/Cx0tDzE+1CuWixxe
MBCBMKiT8mApjCoIvw/DEjw0LSdjSagaTRN0+pxlsFwiy7Q0c+IMRT0GW0reu5SpAVS7yPDLdLk7
HQwuRQ3JMMdBR0upBT84reHWEfWFVWdNUgBAR/Ege8B32sFNZBIGQiso5HerJOO8M7lbGZtb2f7C
4/zKsPyekUC8Fj39DVNgvDw06B+dPSkHBZ0tg8jnbJYwqyPru84aBVw7e8N74PQ6L/72GMlIZf/j
k9gVV6HxbxTGRwfgViqj8E5Fd8BPFrFZpLuWLjAZiSy9U4Q4/VivczFVNPHkVp/x6beUkd8/SjEp
jJ7SYvyidYH8F8LQxCnHkIbDI1xYgvQzJqLEdnjXm+Ox1l+uw7xvGYZqZAB6wqUd/qAqXhUlYRCa
1GArr67EcforxrHvNIJ25FqVtuJb7yzuyZ3rSoMcD9HFBmBVSoI4h+tGQ61sR3RbBfIlmUS3HfJQ
h+z9jxN3wzKYrbzF/llSZG7gbTq2a5oMrzuy+iV1zdwZWh8F42wdd871bor05vc/H0hexit/qJME
dJiDThNLOUXY4z1aMlCCJuQ1u5bQPe+TrR3XWaZVWkpLOf12YevsqFDJE3zxOe9gjEQZIR2mOw+I
+gYHW0HHxOFuWRByMb5bPHr++pyNI2SWQs9vy6YqRFBNZcKubaH1uJ0f/TTYKgmaT61T/VcbnWRb
ekk/7OD904deEuwF4VPHAMNsY94QD5PakcttDQhWdIYvwhhugz3LrPNsW4r3oShQSl9+ysFX24sL
GVTHNTRAqosQ8DpGd4A8xyUI4DwrnQBEz34m82UOlDJN6DBoRGkDBc+9fEaeUJgpFKKkA+41o1VH
j+A4kCwgI3N+DW5NMb0JiEfPwBLFp8K5JTHz8dEDp9Qfo1OWyRjx/Ow1hsWnwPArWViWgAsQJoZd
pGvbPDkFMUHyGGm862u8Jf3FGmXruh0ZQ3cw1ZG8PVLTQGBrU/p0lZq7cC6FNpkWU2NemScz6eVo
koaLGHa2U24tfb4zVodEXoDrkb+yTD+0Y3oVrpN7zuxtiax2avYXIA8mAMKBqjLUyKNRscvE53UG
A3CGV2lQGYk74Efff+uddDk8gXc/gY4eZz+6Jzp0nb1rvbLXJIxRag+oJxkr2Qn69OwuKfljJhRG
CEp4zxwISbpCllkf0h3tBBKgg3OWjF36jCrIixsqUBUNbuJYM2Gqv9dKWqgnlJmBIQRle7S0OuAs
H47ZmiNKXgdTl97M0qkIsDqs4+YnOXl5KQcalxJZtW2ozAZuKtgN8lCYyWjJnmoIWhA55KPlwqXL
A5Qae6BvWGZC7BFJjTWuchYMoiTJ+gdFJD6FqxHjEEtswDt8/DvxeqeG8oE6K839I9v6B07S6qAK
XnZ1eZ8nDjoYEVienlKuau/rKYstt7gvW5CFYbqm7pxydfywbVbdumY3/hpfhWE5w4xHSklSzC6A
VamJNFTan5Eo5Hr1UUvf7aLtLUhiAAnUFNkqXQdf4PGyF3CvjMQz1GOi8x9yV+1dOgxcXCrBygkp
cxjOCu+Y+zqH0022NdaCyqMutjUzzzrW8/M82RU+EM7l8MzSMKe0LYCMkOo/4sR5ygFezuVyTHcY
B7Dh0mgN/lt2QwhKXXGQYV46qlHmDMBN2ECPK/kr+7xOvfl53AM5ZxCxLPpU/zorHJ9Meze/upZA
hNLDa7I8FoK/PoHjyG8NsqwCtjcebu7daKxgyVSnfYWE0c8O12CaEHxPerUiN1Bu1msXajs7MBV9
839bw010KJsH7f0xvAK60xZg6ZjRQcg9QbM6ut9xlnlUiXRGMZOSm7BfJD2FCE9Mfif52lx9mxB2
v7QN/FC3l7cAS4WhdilcjzMStQTwOeBYRQj73vKfamhpO0SoqQvhVGih8PyaSMS4gIbRYabZBtL0
UYia7RfF57sWdxV5X7fAdjV546a6F1Mzol7XdyVfMiB7r/v/iZquQujJ5NKomArxSpYma5l9UU4n
vlzK/tOHda+6KoY9kPxhiEsCOJEA76tCAvVmh1PQfP8j0GiuEN2H2g9IV0Q27QmY6OO9wLD9PypH
2SZq3Zr/J/7pv7RZVimWkgrz4GCKFVg/5Tk70OrigbrhAeQEvNuswCAJx8bTOM/8T7zsLmo0LNuV
z4qxriPY+r68HrOi7nKaQAKIoqLGrtJrQgXwxS+1MFBhmRP8P9xG3be9MSKl5kZ7JUGNrFCE7DUd
OnhJPwRjQCfYEsW09AHPNO3X2iqQJ3wlv4szObCB0SMMFlHejCyQ2xUaityA3t1/TQHdyvBE0E5j
UjHSEvQpQVYQi0uEmme3dZHmYo2GB4Fas73n4PAxGVs2WHVRxt5AJruSbWrTzyYRWkHk0RoGr5bC
4j4hm+Kufe0fBPEfmr2/oeYU2OmZqd1AoBtLHhtE/uUlHtZJQRt9KXfmYYITXFAoJaN7QvSiqUUS
0UW9WEjKEmt2ryn2ptD3BBvBPUwKOtxbVugLKfVvoL3JIZhuU6fQvlfCcnGPHF6s8vwehRtWF1g2
DNkwZrRTQcuXrAFtQl9zTZIRGqkke2f1+Ij7tFAi82mqhztvRh48UrzRcRGLi3N1IkuZPZN2lMCD
e524DDFcVBfFQOANESFKzYJHBueCkwKJFDtTcg28rjG9SXyKHVEnL6Yi3QbosQlbo9B2CFnvuY2x
AuJ/2TgP9QYIgq4U3VG8SNIFrjRFk4ulKHOQyK6HBhdSlODyoSQT4dq9j68oo0U6XCPRgH8pyUNl
w4oHnF9hGE2a95IKI8AzcknXKxMYGttBAH4ybNLjVbnPg+/lI6Nsu94NlTkWz7hJeOdE9/ftXzDM
KqnhkcD2ffZyadvYP7T3vFWT4Qf7o4PmPKe4HZOcICuihYvME3gwEV4AXW4LwxbhSEYBFcHlyIzF
cwfDcbOR+RlKDsw1zBY0pB7vg7BC+zsCGQpcxIAr4wsa1+c0ZyIcnfqiPcwggwrZD5Ss+Fy0ojgX
vm5RJi+B07Lea4+ZyH4/K34jwsgvjDUilXMBYR8EUTkw7c9niDNDE6aUgUr8f/LQT9sCUKbF5/Ki
vL0/+F+s8GNXzkarPl1d5vN7QV6sLSCioWsce8nPqowueglPuxSUIPWCdKhPQLVbzxUoeTPaZzh5
fpUI5mAIaPy5O7Z9B64eY6BZrYe+VQq61CAauBIePAHeUTQ2EPGTiZ6mMJtl7LvrHeu64yiPNdqA
87GIagpsAJEZfxIBX2bZovdvJI3Neqm535lVRTEJZZntwlakh42wA0Js4vlyh7KDVFHGwoBJrz+G
2vBJPO8FUeOR3HLbc3HhHvD3aCYe5JehHprS7TcqCizQISyglXyixwAFkBAyQQNHQqCV/jLDFPSr
+QTedqjipr+4MrYE0nkb0KNYKSmJL3zYloS6cFpQbNYuKMfb9Whmabq1JkPCl7lOCdPoRVkbqzfD
uT1XTtVKaFev+fkApXNsv40z+CRcwrAE/TOCBxUnSjLvu8baHm651UrDXzUpv8S/pRH/IbuGyyZd
jFmp+fhNew2Ze65rRSCmZgE2UhkQDrn1l9BKZmgcMkTQzLXMCM9PE8H/L3n0w85VXh4WA7PY0ilB
yp0ZHqmQP5DiDlL5a/rCAhaZDYW2h/qPgXlZ5o45XlfF+QYFbQZ7IvyVcXk3pMogtUiYPDa2jkSC
2pIvMl0xthrie1zzlkfd7D2/UkbDbq1pIL07Bm9N1DDcSg+Qq2LQ2pdzesW7kXccSNScviiSanve
z74niLCIsZgXKu7O4FoR1FwOJ4/Xyp+M6QMOfGGkBAYKyHbUMudrBtzaGYxg5fv69EuXo09xKeJH
aituXR9VXIVgLdDyDEZru0E5YPVOM0QHHPcME7gSoKmtoUIKJ5SV90FTX0y6lnOR6PUjY9GQLTHb
z6vNNvCpAvKIAx4GPKtdTGjo0cGPvoBs8KmKabwaq5YWvgTGSJz8uLUNMowISLgw9sAdKze+zZvG
o1c5+Sf9WInesJSbMXz0ate6oz9IE+hiK1qRVxPW/a1JyvK/RUy2UWoRnMIAraJ7JLlgjbuzhknj
7NWgih5FmGzvTcEVBzhDbzyJIuFm5yPavQrG3U6Fd3qzbJQWoR/ZbTESGyN5mBRb0BD8KwdpvdaU
5u0buhlFc3oh9/RO9aCg90PRAn81tVFumx9wDRKMchsmvADBqs7rjnDjywXv8YwOX6pUdzX068Ui
nq7dMfGTnrfBXeSTPnrLWmqaO9nBWU7qpK45wHAKXsvjGbI1wIOiTeREK24iDI+V8g1BbxXkUGIf
cyEkOmw0VtR/6+fFX4Wj3v8nVdsMH/nmm/n9GPfA8LuI0pqhbAeSoKltQBdXarqD/jkfU1dw4C4U
AlVos8KJdQoK2Fv1/DyfmNEHzZWYh/FgjuEj4a7xugbMaQBYHnuTKacTkBsf0N0SryTZJzdUuApT
/zu79Yl+gdr7JtwR+RkNWB8T68j1RomHBdk7D9VW0bBL0P6qRgIUl83pc9RqbY3Td632ylOWNuTD
GLHwiHPwizpg5mO2Z7jOUNF4sf43GYj6M3TKdIQV1BFIxflZN3vWqvstdzHaTXX3PSZGjLLAwX7o
/WCxlxRwlsnHiHpTx5ZzlQ7BGE8PAhVoZWt15r7mLKJybIyF8zfhzhAAfGp/aXCBUVeyyHTXboD9
aBxNoV714POMrfnwZNSdqx3ev0SCg0DBR6IbuuJKaDU4XhK3oIDXZYwnHpowmQQ3pfAjAIcyaEx1
HVOimEeqxCnE7zAYyBROo2Bs63Wj+7UP8Vd42u6+QV9HKT/d4NJfti/W3viBMshejmI4u4gGIIyA
GnadE7fmPJpx6A7rIhC0QW5mnpdYIfVmjUuBofagw4oMU8z0ecmEWGp5agWMUYXkqtppIn/I67yv
9J0V9jqxLUqH5zXtUGtTSuJnl7+TVKjsBE7LXJFRRvz7Ut+Y56p8AkjKqIFxvCNzfpCpiw5/PO6i
cRAZLVFzpoojHK8I4m27rzHbZ/PNuWsjwnyMXXaFJjrbyBEsUryoNwaWxatGxoNSi3/xoQcbtpil
fATzLSNxZKxBSG1mjym/a1AAchc+t3cG6Jq6cKxngVfdNRLypfYGcs6q8vGXYsKiijlxmazmW5P7
17GC0FHC5AsrjjDOozeH/z2cq8HzQKfkNnWPn8naOvL52l3XY3BW9RQ61oPtXQYUa0GEgGUXRlOh
jzUPI+EkkUNElFPy2Mczc9N6K8B+qhThZOJoWoaqcBfReQn47bKepo3w3Hr2c2rxJsTUp3nF1Uax
CS7XmSiHjG5g+ZQ+q3wOfx8AvgTxfGafnvzmIUQ0acnn4l1s+NGJ2l7IZSC0vKdraM2EC9/3shqm
YE4w4hw1523k9NjH6zex+xk8reTcf0oUeA3IIfBzCFwiLDyMxtleeHeyA9AXrwpgNqVFYgz0Z5rq
99vY+/jd1WZ/HGHMSsmpIR/udr++BI3nQ5RiQRoDmGyverpD8efe4hYO0hNS5ZxWBOAJ66yFDVGb
qXcY0Y7CQzTWtHkfAK3lwq+xSanJi9HuDbTFzKqjVv5PCJbI5W1guz5XQzQ86Y6KzcZNKlk7LTLR
r5I/zDojeQ/7FFOeDGpExkXTXOeWM2Ye5IcwnEsyjL9PEGCI1XTFvtKW+mzMsYKQX9Dp/+/oJ6v+
uXWvLZfJOXUTDP3qSepEhQofwl+KSrt7TpxpWYBf9X97MXA7OXbxQ8PmT/e2RsMhgy+GIcDrIl6D
Brfqdj33/Hn2uA790By7rFOVuo8VRK24zAqXGB1uyq6NEESl7aHRdXbH3qHWyRowmdSHfZxqVMaA
y9hauHkBR89LrOBgBD9fh7E9Hbu197rylAaatCoyQ2lZl4ADeJcDLi9UGIH+AdWuLIZVe7rlbk8U
0wfBc0auyDw++sUrRgtcZO+FM8HlRw6l6PCt6HEsb6elCv8CpHPKmJR0iB6Exdn34gU5x1OVBuAz
8AEfvZpDqrE2WVOA1KLqAXfbJ1HdjgcCO5VJKwxS/pugDTIysex4F+lKfBKbO0IOZXa3rw3A+Y5D
rOp+oGEyjOneNpoV62/WtBvFBirklohfvDELotAq+9MF+A4kW+6dgkGuUP7gX7cRP85jAznNIJuW
5ee1UOZmVAZSiBqwt/ap4sqJC4IhV6bhPF0jOWCWe/d/axALwBCinzOV6rqn7rldOdFd5XVFBf3h
s7FiJrmXKK19/kKfc9c3hKyt/YupPe4vQ300cjwZW1vvOtLKMBz0LK5bvbxwuDPvbZg439JweAPL
VfqpzeEyS+I3Dhlc8eAFrpVxv3ctGRhsjX7voVjrkoMb5qoCzmPTyUU+T3QGfJ7/shXOS2zpBAJ5
AzYj8KmcO/34cjOftWtmW8SywfmdBMuCKISbYJuCzXJhOetYjW1l6bFjrojh29BRrk/sQm3Uwoc+
rRJzmeBlgaer0A9ZApnHprkSDrghtpUgwCJzFBhpT8Mw8e2dMFMWmTvGTMQSMB9zGnODXUG/pm/w
Wfdh7wc0qoUG/itmJOqK4y21vXHRjHgTkoqSHbDB2NT9p0p4hZulmqBDV0aCQTz+h8+6yTKi0wMH
56zm6ayph9JcmAql4mArDMFhz0zPQMzm3CLLGXeCYgx5X93kwn5rtEfdyFp2yXlsN19nkltSbuSU
OqFpxHBCPioq6X660i/Ob8lcgUVwjDqbppxVSPpB1Hjh66thl8u9Ta+GTJM+hFlparcMuxN5Qf50
n8zeFOfQ3mGiFUW49NgeNZVne4osDFFHF4CiR9bgY7D48ZWhiWs19cgCBlbQckW1Kicw0A0ckLpY
+2PVFBBwC+cf3rkly0PJqW51+hyptbwNdcbtGHcXp76nigkVnZ7V3HNF0xxmuYtntwff3zn4PhvA
/f4pOWCfiuDsy1CLSC6wleIdxn83Cr9p9BrdQTxaQHyc1Uo0ebaYDeSwzSi5O7D3sP3uEw9FgaSN
l46UgoZXAxOHzaLhvy8zDwDr7wAMo6Dp9yeHo8ktOZswaSvUasZaJ8SUhx0HXg0nQv+Ls+pONZFO
lxqkTdA8CJL6rucC2nuxwyVhztlsHq22lwhMqv8GeOnYtPBk0mXno2i/7l+PNi80BuDbbhLYLlPV
MkixcGmAtVDQlCNJQtB4TW04YkuHHBu23q/DXdjmvzaeCKrd9croI3HiIEc/xLCoSciyV5Pxdms3
47ZeN3kjN5Xst9KRD5VG7tcV1/sTkmnzA7L9qpmVZhkKxVFGpMBruh0uBSHukUkVNCphuL4fyq4j
GHn5Xt5rttjcv0DYO+3TdOlo/HQN9fOyxT4BP2d9hHp+Cj5VLYe8E/4VQ3nsDlgqSd8TD6cKGvAH
kECT1cjzZXVlvoBK99YaAccFbi9KOx3t+5KoyQnV92MJ3bB0LtvH7HBLQlOn6kelH+f2MXDlgwfY
C3K3HDKZtyoBmWrbhe0+nUe3mn0+3gx8k4nezWUFH4QUS6ElQw/NIVKDurJNtD9ftn9d0Qs2XrGT
HC8nhmj7WLTBBKRPpdaWkl08pOMX6+lsfAjdMQpn76IVAo2w2sDok1Ts8qEU5bAOHpIixU/KAltU
lzRDm+Az0plcGah7ECky60PlJC0tp/kTQj7SnRc2dOO+XrLbO1gyB4IZyrNmIsTNUp5ySl10d4TX
bCQaDGxlE5fjKmOiKrWHuOATTCWy3JZEiJKwDxwGfZChkx03mnXk8ArOejrTC1zr0Y/4zsqYRokd
+0B8ePOHbfpNcfsWrNNRgGSpjHsZtqtOVRrat5zwJ0i9Al4gT5zK7neS54Dgqnvjr6BTT9MUdJ/M
bPodMfh8WzHlPRvBLxD3kgX0clF+pFMgirIKH8ZzAcgv8XOV20bPp1zuVBa4ggbuznF7hBko+Mba
WpW08oVjPql8CHZkQhQLEECNMoD7GNlmEhXSxkZvMqK7XagQ43LTFhiz5s5nPg2mRFugnToupqYl
5+UzOB3t6RyEpTc3tikyDTCMI3QtdNpVB/+R5Ws5agxLzKioH9ZbnnSN9X9q9EDcWGqjkfX0RqHV
2BZK4Of2Q3ubG5ksmBLPyu0RWWtzgQ6lVvExBHqTgPYHj+P9aw8gALSbsUby8Vk4q/1dNNUQJI7x
CYezpFYCo/OXuHCdEqApai+e7djVJuG+rU+/0uMIABCeZ1V6CP0DOZo4mXo97jBbJR132SJnECbl
zQ55xCgSUTEk1CjGi2wNAr/i1nZVCq8vBPlHtCcfjuQIGyls7ZwGzXneSoPlIdD9+xQmOyp5MHgA
zSsEVTP1EfX0il2DUN7oYaZsEgulQcj8Q5o4e+KH93Jy5Ook9H6V2V4J16ujU90t2fNVjLC7Tx6r
93Uq1j171XlM+v5I2q1/xVue+7uDzijQvCIGgalNXQFEeDq9qJuZl2xGlafsqpb2iU391KqGdYeg
tgjS2S+3WzAn9tQLnebhNCQn7Mj9eYw5GGI4YIVxSGXOeE0EQHKG1H4qJhc9urkQwqqdxJje3unc
PnoNt+1QY3Bdp1csVYjsi+I6WBQebhoI4nm8a/ocxCgHZFkHqwqRbuocxAJJncBmF6pBny+w0B2M
XZprgoM/mq9AxiCQ9Geh88O6p9n/k1AB5wZ22bHoHDznDjfjzlPFucBLL0nUiYAW8L7pS4KUMVQ4
bYMIKDOTp4O1m4pQLcws6zZWWJERy7HuG3+giQmCzDPvaUdrUVcE3ABLV6OQMKZGER7vpQwbr0BV
qpDXk+Y627GbuFgMbnfdO5WmVdO0ruil6fl2NDd9mltGZub1PMjMAiEy6k6sRZZ6AA50J2UAe6eN
rhGF1uwOzcCOKNFB5JlMroXq0+mPBaSQzBQvRqmDIXYHqV5pNV9T7Ka8Hjkl7BCWFUlBFstn98xW
mJy4GVpU2En0ahLB6yGIWlCvLpWLloXYhOlKWtZ79MrjqxDLvZgMfiXBDCk70Z3/YtQ2Rv1V4oJE
Rowki+fkk+XUM6fFWqJlBgtGHWUnElEqynaVbx4b97hxJgBL97lM+28v8dd6DFVugEKYQUy6QtZi
QWMDBVD7VUsNnQFjrJ0aKYveYUDeuZloKsVQL7PZL+/3n0fnREYT9Vfjmkmex7lXteaEXL4RivrN
reMaKKIgnlGKJVjHhFA9316WWt+eYqAlH+PtguVf05qTCe5XgE9AnImXr+/Bhk6rZtISkYSBbC6N
a3jLzbvHCTPCPnSymYk4qwGgd9i7P4cIrSNztX+1GW8thGP/K7462mxTrodCROXFKOx/FI9Sbtit
lcRU2InUt69UkTbXKZ7KP23vh14sJYlAPqeSxsidKq3S9EcM+DRi4IuKbqfhY2ONI0ASDobanalO
yrXdFg9pI1afHTxH2VrVbtoltkHgMx67JnzoOsuPqQbqnnQ3yPGHo2IdkFSeIm00WQisKugWYYTC
4nE8gLipFyN7EEJOlz585/jlXDZXQZgZSLcOd/II+BQqKkV6HFlwOZWsHKSSnKkjeKYM4/FHKPC8
frfK5VEfhEQ0WdLykLze7jCk6o7MkjUNxrBXbFFdRjujXJgepKkXIjoua4+sqSkj8PYI1JHd3Zgq
CWZKo/IuK/58WGWC1TJ/XtUf7giiTwffN2Waxs+WkOU7ZtEWDnzv9dHVSDOOenNFdv3rBCu7Glf9
94DJfOynzXV6yc1iLPj0sq9Kr2UVMPG6Nb4NdLBqZZhoA9l6jhul3ooeK+gSDWZyI4jX343m4V1r
wgzue/xpu3xlazJXObiPwe8s0TWW5+zoX0t62tzrnxwuNqDuJN2hmFCdnwXU/PSNn/1KlgzwDtOw
ieFGpLo50NLwqUuAAcGczBs9aBNZSlXlj3UgPrqONjzjiMN7a5YbTWmph0SrRsGQZbNQvb5lYQpE
k6xo+cnfvWkb9qIQIxQBBQIyFiDEYU4GugXU77SnKGzbKZ9XEELPjMEpgxdMD64NibE+yjLZYeEK
+OZxWsyb0RsGFeKT4uQrpe/uCBaA8j+AYjcSIRAxIUQt2LD3L/Lwl+5NLRZ97AncvJ4J8KersX0C
a4mIw+4SjVm01jGy+X8+3X52RS7kLckxOFnYY2p0JWsrd5k1Zhh94QOd/fBECdUEDJ5McCjKw1ot
N85u9094QFhzFEXga6P4Me9FkEuXZOnl1LBMehZ58KvScyKtuZZGOrQ1kkthqEWGMOxhwLH7ayAG
8uOD9gLtascUNH4XyLULKxE/IQbeKvdZBOj1HaxWOqs0siTsJFm/XlIY8yFSriBHR5RwgeXoJl1Q
RxWsAmjf6FGVaNaiRdBTKurJpsPaP1nUYwpTVzgUyhC6mOINBcQUZzI+JCE/uY3zZ2czuDCNuW5Q
JW+If+6bNYu9073EntzM0Q2CAuUTMYYnCKoJihWpP8ORXQ7sfRHoGqP6W6qYjDeUk2yz9uUqsfoy
n0hsb5otipkU9Mwm0INre6Y4s3XEV2gs6WKGlVfSAd0frgbFBP6AVEkMesg7L3axr2RiZhtHZ/6d
CagOGetM5LJ60bCz8ytelwx0KJYHpxQvGymlj49B7y4kCOzVCSTDgqaZTF2uSjjsv6TGjhMWCGkr
qfVL1REufbyaxm3cn4Q+6ax8hjMnzSPeQT8ie2P60ky4kNqRc+jyZTmozY9DDTC4DpPC4F7cY9Sp
1/EBpgSRqlMoqI282g92X8brNOxhfFwlNYM9NQlcY+/ORfnn5YhXXINs2U4CLI4kS+NTihxY9hBc
UEhqXTrjP4KK4mAsJeDBTlka+yiu6nD2ZHOhQVmu9z51VNsn2+7AHjJswpHIScZI9ayuXf6/JeFy
IsDOWLWt04Mifkym4mwUyQVe8skFCnTAv6s32sb6xoriIlVJC+PS8TKca2nV1Fmc0diALXy4il3Q
NKbKe7KTZKr6ZEQHkEXIemrVZWc/94HzJg2DIbD8RgyY7fYPgX0D24IjyRpPwcZtYQxGWIaL/O+z
82PWjQAnGmhev7tXNiky1manLxZ54Ajsz3207OZsEThFiV1/TyP0keEoCsCNihlssWEIur3qLa50
NItVQKkbC+agoLOe2EBP010qi4PBJHjh9TW/dJm9lo/IYl4iz24FNvAnY/zwygOP9kyjtJ1PsbfZ
gPTGXfZri8581s3vLTucRkrmnb7IneN6BcV76APhtPjbKXfZ2QIj8lxCqT+lUV00sDNqRyPqiEVE
oaTSmSJGwh3sDAomB1Me/laJIogkubYxOJRoC5MCPqb9HA6vFpwRFG6nzImRLaCXV6kSXdoRKQMP
dleT9+biVKSKyU2KRV7gmeoaaGpVJmGR39pNNwf3F/OwH9lyYzWoPVwEm/2iLFV7XVhbp6oDK7KU
CIcl6hSD+JQAjQryK8uDMrbfhb8G6jtL2LKF7RFaQSMtNBw6z6cz/GyU8KLlFyooPL8aAuV2fBY3
a6zn/5Rq2ZXYJxekqrg0K9lr9gsXRe37TD3QQQD41HId0uCOYc3tB74z7a/wtNV8sDguGAX8uHrw
ovL/af8WgURRddxw5IL2fR9ptiJPXKzelatgC0HNQOm5HqQ833wCDK2B8AUXyfjOtgQnmtvnT4Jn
P0yb9dxpFEVE3Yxk+SNYJwsgTT5cbqoq5mRrALMNWClqzkCv1Y0ztPbFBJwczockUKckCf0+mWc7
v1nfe9JhbOEguyuVmZFq9Ij/m/J+fuudb4ThuErXtuxiQd9ISSuL7oyk0VYhIXfRik6jV4kEz1ro
eIqQFTkCsEcKd4p72578QV2RCNHIx6pQ7NokiAWbv+/dmGzyfek44dSdklQLc12+uuKJ2kxuTJEC
wj30wKbNto7ICh9R9gOW/G6gxR4pGZeCGNuvui4m+IA/1/TusJPS6GGXgYPcO3jfsahbKvFDO5Wi
vE6B0x60lku2maHtTmnvlt7KZE/qB3PUvRFz33RVF3sEKzucQw4uAW0Is4H+TOuNfG1FRyZHcmUL
PyNKgKCjMj7DVRLBGJwkLn09ovNpD5HldF+Cif393zsy3jl0f1gL/5Eu90ZnJzNJbkJFFRbvph/7
lMoZBrz4fRHeuf+hatVsH5hPJnHCJUIknItASnZw69T2BlGimEz7ajNdW+lZPuxJyFHjwV4faHIh
PhuVkLi+gBVyeW+XU57R0nsDyW5b5YAnzzOhHlx3WsBSNd5yM8JNpVj2Ns/wm4MUGuTWI22dNErh
3wROQSkVK5+a+KRfeLOeubBk/V0Wk8NPRglwhNnS643JdtkbAjNEQcTHtu/9u5mMkE3CBkYTMfwY
bQs+lM5Xmc9hhVrqtT3i8PcGedl4yKSIA9yKpd621vvefXzNgCE95fichglSQGnN70xRQ0B/RIV3
QR2Npeoamy9BmHivZ50PVmDm/4Y65v7FjjDrqfmkD2+TO0YcRoc6HEfw1Aw0W470GsupDFU2lMtd
xUNXmMNFy3AATNSzoxyl2fxljcRrIzkn3zy2EFf2Qnf/iZFMp+5U5J5MHOEzP1geE0jZ3lKJoNWH
ieuZShtxZ47bTh9dxmoSCo+ajSbklAGJZvATg5bpz41iNykH0EKcq89080NusHN2YFzb0GZ9rCrU
gp+7rfzGIqp5yGuVQYqVn1WVsAWdktOT0iEcKCYT+emXRnK51IWXZrtAOG+4//FTxwKOaMXOViEj
wDiv6f+/A66ezK2ED9KUImPYyFMXos8fHuQ2vxqYPeR0uNK/scBYdNVHBa37+VQNfQxvZPBD8JDm
gM8v3btZeimvZeXBMe9GpycrW4UBUHHJAYGoIwqGoGkDQ35Ot235Iel1vnnsYhS6qWssqOvdlUlJ
2HpMQyJ7mCtmrKVwvwlYPpbnv2sF3JwK6PdgdJZ2gPTDkEWV+UGQ2kOLJOTyl6bYanu4kF2Q/VLr
T01CA4UWucD6zJJsjailR3fcbvkbdnzs/vtd/CrA1TckojNHRq3xp6OeQr1lQGNwe3XYdk3apvVm
tnBFMTn0/QuIsBFI30zf/I8u2N627g3SkHZpSQSMt3lcrwxN7sL0k37uc66J5d0h29gnf4hcr1H2
w3aHQcu5lyclVN8Zbp0GsXJyd/gZ6KP2AKgqfHNQE3wnfFgEuLERM23VtdpB6FeMfs3V15o1HO12
QIWNA9EvkibIQ5vW0HF44y7+sUP+GtKK8V33nOv7AA1hqsdIvm83/Otlo07vutbCxgdJHe+JeBvV
L3pUOSWTgBFlk+a/BV2X7p6rVDkPwoXerS2Uq9bnB3ubu2YhVj/6QskIgr7YjlGjOqSg8jYnBAo6
0XjeIp+8K04YTdbhW4xkuQ9QfDtS0k3anYXWq+zvs4QD0LpB6O8KtsddwUlBmEIWLS0mGHuTQlIA
eZ8UQFRmgZDT/VWd7hazxM+cn4HNzzarGRrc/tgNz405v0tKntopZ3cTtF/ymharBkiNh14cEXNI
krfaA7ueQ5J2edE/j+kwSiBQ/XY0vj3HA/E+HlwWmMd+Xr0e/TX+AWcvJ1PNinL695ApTXyFBTPD
zkyThJNdWwbA8VO6SnapsZOPIhvjGJqRS12CFJ9n8mwPbh1ybeCBw75qcMpNE82VPbwCh7IDSkWV
Hr7NtYVzBXT4JfFUYMmjU7GIFykWzbZV8rlP8NZqfEfmCFEt5zmroUAk7vwQ4TCX9GsBCVv/9oPf
xjHk1CBkUqoxi6Id0rGAumuwTfhL4CPRG0iLUmdnq1ATDJL3QuINHvZH07n1/T8LQvyKyd4W6gYB
lzpokomMIy32rPkmCIFw98QD/GSZL9ydtBRNa2AwhbLEsgMr8mlEKT318DGsM4wXxEtn6Euh2S4m
wYoLFFDKxjiOP8ZcHOgtGNOBK70xynUk69wS3R7aYBEd4CiC2QbKK+qpa+Z4OUOuHof3FzPCbiO9
l39K2yAAC+/T6FQmk0v/V8/pEK0S+T/FAsEIVxSqvIdCqK9e/abK0C6uQ+MEhfHsE/ShyKJo1vNq
uL/otohgFl/HgVqkNvSTEv4vtTFDO6NzifdETEXonq89rTWysgHajoY1UkNzr1BTGzCm+QpYeEau
ADWYQJAgbw8XHDN1prRtOOaMkWqKtJTXB1obHhYaQ637wtr+vcwjKdNsaAGOqWdchahjg2Vcub9h
baFNBDRwf+64d4JY7lECcZaoRr7g59fGIVmXZH+kxbxC2zBI2abzjrffa9YCfhxQP8knMeDRivR5
7Y06uXi/FN/TWIoZ+e3/yEHx68EWw4q2t4ESSVMzHhWvyPmxjsMtPeZD9Nu2uAqEWzw16ZK8PZ8l
UDOjM5KCIMsnu+9uflsyYIvAgCQWcxAv5Q2XvjJplRqxR0QpBExwKHGHIDrBkBatN/sBN8Z9Kdyl
AUUWdsb/nZAK0w0x6qAoehjncvX4l0YymT7Y+rJifSjl/yJOnkDbFV/RpIWiyX/BgjF7DmEIUB7o
atjqJPX0/EzpdbaaGyG6HkrwHqwt8Z+h1Ui4eQw+7qX2oz6EK/sGjscmedVX1k9kHeMzewjapBMM
Z0Gw8j2B8byxlatdGC+pVbTBEAGlnVB5qyhHiKafJNJjA/fuMZSuB2qYs0vtdwiKdv3HBpDrZYYH
98ictprk2nV4yBSkXRsa5Ar6WTzKOWGx88KZs7alKCtt36+svIznaPAornxTatLEpwLgruNLB+qE
nymFE3aKMSC+ot5GHpHAY1jMBblObSMjZveW+pvZLLq3wGevxwYltg4IY0tjku1StZ9I30V9z2h0
An52XZN4LAa/EKTHvTVBM/Qfj8oDFWY/wtdL2AWQclv/Ufpb2/tF3x/G17Vy0720fUY2p8qPPaJq
4eV7of5E5zwHqe03E2Rgob9ijpu+NEJwH5AroRDDPtrMvReBIs6EoDTsV2MNpn3B4onAHvOMPPTa
aG7e/5BnXP7v/x31WXoqBx7x9B4L8VH/dTwhBKtVk/NHuW93J6Qwpeht5ogfp2DZWP3kWG965Ed9
eVpRF7DXP7h68Kk4mVK02GyDILoyQqhnneN/gTw8vYtp2reE3UJAEhyuHuYWD37hGyLf3rBxAXLo
Rl06yPcKIx66vyaRYrPlnfUHqC0CP0R6Aunmz1cMVtWmU8wfC2RSnPlxtlC1426h5LLWEpnP0VZH
79M36LvVcwFbfS6Xksoziso1ipJ8uu+Gs5MGbIiiXG+g7GTL3Oglit+/vhY53taM4w8bgE/CsOXg
wwPq4p9BoT+Z+mKihUw4hr0oE5r9r51uCKv3P1VR3V3Z3ivOXZvyZLAfatQKfdKDshxqykLcgMEy
Diw6tLiOMS11B3KLt+0Z24ALjGcLiUPzHPlZXTvzBJrmDYiCAdB7UQYjBunbaczZKZa4OUc93VtN
LKF9Z0rc/ItHFTYxKtHO3aVqHJzUVn1hnXq/DAPe7hloLYKq0n0ekcPGZGpV0vTfhIJJeFM42nNX
FyBGnthsq8Dp98cHgxMjPKFPO7kgfHJeoGMzaEVDxkbuKVqWDn4q39xRnfJeFMkNjuSV3P4+whCT
bilqPYaO3Uv9A30PWnDABpzH9gQzd38cbgYBbPxJEWlm9xe1b8NtKebUPd0eQt45qs+lUGIMRI2X
+Zca/2tZAf2pTrC2+BrnNqKumM7KbSA1Cvovz/JVmfbfHhLsPorNmCJ4+HZnFeXGWsSbfN7lRM1G
uh7TepfGxeiIl28PI/42sbr6448XLe/F+YNan4MFYfHJfYoRWuo7qgyBOKWo4f/NLX1XhcAW+oE2
qOR8Y0zDKexgKh7mXxsQuIF//9MM4fnBKzobn8cUfxp155fEJXcTNNyzvEc1myKfHEfA5bfK5MdF
ZO8sBKiw4YN+FM3se+oW8CnkR4ew6cEhClWf7R3ak3azbKNzSDnwycb5fhHbif6Udkvgco1ZU+hf
yyXKfw2WUPt0DcDcJ4n7kJaiA1eIlJVyqyJh23V/kpMx0XOuQcqnWUxEWhRmQX0qlWowBmbreXhr
VYNP2fLP5fRdYe/SE4AANAF3v+ylHQVmzxuj1+noZx3aV1Fz4EWbNVnpUWTHwP+nzlc2CXf+Ss6f
cdQosa0C9mKVcdCXStvfl6lkUrspz+fscK79Of/0Q3MKg7gTTQwSVZFgW2wPCZ0ZRqNGjyFD63Sv
VQ3q39FfNTckaLzPjmJpQyWpeKFKUMWnQbfrSphMDDtazqu2wRm/GKnaISVQ6X+M/bbip+rBA3AH
XdyNDjT+nJ9N/5GsTMQlzs9Nsn5breHJ9S+kDGoCsfCtQtgQNW1GLjuWQ/oJ4by7j7KwSmEvfyGL
aApUeGKcTe++Uw8lHqDgqPU6uM19xiDAoOHFMckkXPjSnN/JmS3F88jmNI4mTTJzaO8OAOgQaq/A
2mkl9GtU7dA08u+jtPSE6pFckPc3hJo6IBYoYStSvBY1geE5+Qgf8ZTGTpbfY8nVwquxCG6CHOsB
s4dcQj9OAw9Ug5A3eu+5hu/4ckRn+xQBoOhwNUVcYBBfDcDPM/k96PQvhAzCGqHJZ25xCRTMNtow
NX7sZWx0XTT0aMbPPwpgXLn9g3FdECFdLWnjRcVmSYrIeQfeuBJfyq7eOx3sqeQsusqhl2jf077a
1PcYSJGS1b4LLiGSwIp27FiZV9R4P2YuiLNv48w+s/o4jrJfkMC5YDYzwnQeLbxRJJclXqexDe26
6Gv5JGSCzTZEkRls4MRmir9rM5s26psi5eH9hSwhRliNNiEvfP1YFYEBsOaKkJJYPCAOtlQpUUam
nFBcY3rf/2JERdySrtCxcp/HPRlD4JryuDZNGAFqmwz0iDW9Mk/oo1JIIrS3mNcPexgvAvzy1DAW
ozl8tftWaODq7kwUd2jqFGRmBDAMKASkiPCWOlvdjJpSSuXPyJU0oqamEaWlQIyewD5heLEXUF2+
A/ck7OM/KfVuU25neIqZA36uX8b6/tlPF4CREnBClrb+j0K3tQZ1Y26F7+hHaOEL1Ta/TXRYPUti
7Qx7SxT5C5UybVo7YotwbGnwUVCDA998dIFWMu/IHYKyhG3a5tZqTr00uTXfkIRsrhdKHDoO2tVF
h+D3AHNvirw5+IbnlLBkskl2EFzieSeq8vlmS2XeuAP5lG5vt++SUBpogGWYp64NjHQylbV8k2Ie
QVSr3If3x9e9nJoMSr9VqGMqoy8zM/yvo0nTzWEcv7ftaXU0mEaWzTNs/kZzObJptm4AIixLAhDi
rkL/zB+L56XjoF8Ci4A9jNrOeZ7myvWRcaO3K48pAbX/jhbjpCQyZPQsrpV8uO4H116D/bP+ZsDQ
sEnMus7B4hWXtTlBFO3aekkeLp2uWQs/4hLFZfu0v22zu7UbmUt3fTN0F9cAodfB8+ryGN82usH3
YLPumtGdd15I10YoE8FeRfFjPLZtFmkgGw7kp7ziBiXnaqWeNskgjNhvOwFiRzsfvXqTcmAfpbvF
30DwoXoRgcFEYAd07Jb7iA56ySoSTr/LAxoYUqNXdL5GDLCmFJP9k9gUFlGIPU5+gzZ7ysIYKDS5
BivEVgg8wm6X7xIgK+4UnWx8Any1MZBUVgPb5llLFbcNBzl4Glkk6gjMqhKQA9Fc4OjSR/nDCRh+
BqJHqhdOShbiBh+TZLbJ+87SrAzqAjFVR2ufgMa4uFOVGabkjG0BmFOecL2eRfG2mYF6H+inYh/v
UGQnpfPyZOH5uAqxhAKA2WYiRJ6Jmsg2/GVJJ48+TFS//fKLaW+V6BsX1GvFsfrT7Of7zwjsVVZ8
pQDOfldK2Aga5oMyxzJg+23DiVI/gH9PdLn8QQXe5yFNK6UTmBlV1n4LtzDC9vZRXfx7ihfzFpqz
fiyYWuJvo6rlutOh5KyI/w3jlN+RNGC9/0+atKVShDQYFe4wbxJvo7Ea3c4nxjCbeEGF0RBEz/vT
Jia2MzCYy9761fhaGUOwTA7V9pHbdEjWFdBJ96CnUkOo5YmDllCE/xwmpHgjulxdCO1h7cdlZKT0
esVqhMr2ra6lyfpj9rA9vDzX1pIhYA5IwsYNtLcy5DttehtKvxTfHZjK+eToQmzhnWxmJ2HA7n5+
gj+6L3T3tpeU51mcj9YKgjAhgjuoG5XWIysEswkjCM+X+Aar0HxHN4np2IdhnbW0eXfy/J2rZboJ
dwyjWFM4MfK24ngWmOXy+AB9Ns7cJfkEcriMSfw1RrKINY4I0tIPPtB0juWiexg+1432jwdsoPYo
s91shBDbpGAy4tYIVl++dTiKg+d9FizlZdGNSLUzWKRHxKEL/hMOLckwqxsvf3hbocuQEchlBruX
0kfhP6Bk+1hz8AXYDjXWcJIbN6P9V75YAekbpYKJEhufCKkMlbeC167jLSg4QYrMkFviEwwPu28X
Je9rMrBvTOMu1Ol76nn7y0gnKkBfnZkkXtJN1BuJX/YqPtwcqxMpMbFiRhJJ25yox7JDm1Z9Dxfl
tJvpS9YHn8cghEJ+9l11KVTHfeG8l0MTJvOhoIoG5vzzKnV0WYKm5wLY45OHJluY8o4+y8dH2t1q
TkNFt68Ial+YFz30t4Z5+lEDOjon49UCBQqU9gN7Yb9RTyv96nDJ5Ow84l7mgt+h1P5F0LNwU/NP
ApWPZBCrucDcitmzl8lza6pIAvI/n7ONyt3RbRcDfwhJXjx8Vkw+L0gqDNKVlchexECI4yqVxhrW
Z/ASRN86yNmcZa15VXeUl5RgS1a58UybrH/UiSZ2/AIz2ts1LjpWwo/yM8h3UldNz6mcfiMYS+mg
ZiHVPPbqNpkDoijeX77rZ1/SGO/4NdJ+8D481U5amccCCzsThCgY0k8/b7tAmUFMbTlv6apI5p1T
yOC2tKwRljf2p59I0WzlnCB9QjA/CE/BiYERJkE2ZrYDA7j+/fQfNz8dTu3P2wT0Q0DfGCyn3f9r
EAcwzKzfl1k4VpcDjs/at2AIT9SjpGcx+7Wzl9VIK7Pcq+yufdznF5X+sU2obmE7tMyTzd2FSLkx
QeWq30cGto/M3y1EdAwGNoKPSeQyVxzmTuWgf1dnaS4hgtWrFBr5p595naieXEdyHuk8Cw+ZJK52
+aN8KTtkhKfl1pE+PrdBX5aotV66y4YQyDrgetH4N6+c72M03sAT216LEp+M3uZoIB6mUgkPrjwN
heXNEnxaWF7gJCLr3v5QS4RQLrdfT2NZQeWXvLmwtDJwM2TifH9yuOjH3IHQ2y8GCXXfPPYslwNv
5JlZsRNx578LwDmPFNtdBhPsJfEZZpYWVBxJUJM52CMOWM0nlWkql2WdYwVL6K0/JfM+PqCR5fFZ
DNBJ3zYnLUUJMNEaSz/sW+NnWyfbIqHdlQQqBPBVy4F4j2o/Q+/MKzzyFU5Mu4XxNklu6C+MEeO2
nt1Z5wbi5l+9hmcYOfLwfH7Nir0X8gAr/7lzRWg4vkDX2QBpc/pADNEppt9A0uWKQiGYKLzDpGhl
BosoGLfnV7JBIc06ZcAbGkdlnvMmEeqtsOKVVDC9NHSkqvPBzhcx0YMzQRtRRpgi1BIZnS+dJCOq
vC65azZX5Axbr6NkIULrrXZJQ4lNloOS3w8ltTM2AKUKbNP+J6uGcE3Mj6ihuk+wU6fguFWdWrlt
zte8cFHtYZVYK9VVP9WAaE0UmhsZuONxd572S8PbgBTQ1bOPY6TnVSNStWCHymZB61wJE1iAsuys
e+6poL7591Aaln1hErgK6aj0BeWnm24cEw4RpWSH6A/jCMteH5u8zcQxXUg7RwN0dGpS/P+xifJY
ScesfKU/FFeYAwOQ2ddgmPMRMoWyWwMnOdQA/MKNRPlbwVk8QfoNOJWJQCHzXRt9m4NSaiTjP+Ls
QF2ChLNpMx5F/qz2mhPMVpDbhOXQOlU7ya2AcR2oOn6rYvExSPzkBL1USoW65HEeSbO20niL/6hS
tP7oVyiJgAThB2mzYeY83DVp2KGJeg6Az+GuSywt9w5ErvlgaKQYSidx8WmcaNaKLnYgqhuRaxLB
T/5L+jYvfggmsQgnvxoza8iqLlH1mDLPB7FbRSyVmDQFgbtZKrcMsRAYRqo6Ro/MTwbOnqunn/69
bhbv2ZES8yrsIzAQt84XKI6mBd5GwFD6rnmkzgMt69t3J7p/bsxhYiNgnsABxsUzCAFpxnN1t4AS
KEQ3tzSVopCRdXOIEBWaDI92Sz8/nTtG37ls2gghziXNO7i6qZGqErBaI3BhyLbR9S+Fs4mxir6w
5UkeEK3PblpyDFm2JeK8ZYCSF0uoKtSA02RNENgbNtzNMiPcWjMsdw5qyUyGrAXWad5eoKFc5Z5K
LzVjBR4RaCD1GaEUlw1P4xiYK3FbQf3qifk1EUupF0rYUxUw5sXSqnq7xbwPhWfJSwd43N4WGdPC
r9/8n0Hwu//3T2r398VdOCHHKjKaTFnSszFY6Ovx6hw6XgUK2bGeUMKDGXXujA5aSujhJtuPyoQ3
9unafV3N1L0aZjF7q8dSMIjbwaxUP+qlU51vbIDKixgtxV7xckvogcgN9f7t7ZmbOxesjyU1xaqe
hIwiEK2rKyxuTudP1kWQDvZQLnYllL65hHl5yVl4ZVVDVbDRqBUrrOjKHv+EfMFIvTvpn3JXYjGk
3SPD40hAe17UWtxIp9ysdGfkkN/tEbD2lXMhiFhj6KEs0fzm/nIwE//MmTDL8v7q57A+JN69oTHm
GEvcXgsO9diMJzOQ4yVPpOlQGSEar9eaxReBBlffFq8zs9lzJh5ofoyySE8yTmdYZyDXA9jY5Eq8
7mtq51p1ZX3zRvQnYfzO40YGy1guMHcB+XSc5BYJMNo7YCjoeXeQmAN1mhpbrMucVQBXP0GscsJu
9n5kibRXs9RXgx1nnYT4A0YUNt3MNfiY3Tqv6NoRYNeTsQGtE4I1kBF4w/XsLSMr0bPf2Y7Oy7kB
SeRDSgtReQynL1xpTyQtdrQpEEpfhbzBcklgtFdxdby98XHy9eaRiG/Fwq8d29KfXdgkssLzWnLg
CJPy7S7xFLumbbPgL6NGRamP6O5w6/ySl5/wydc7l3uZ8AWP6I6o7hLbUjtbyJYIWllLe81SGQJx
XKKamNpFcO4wqq3WDtkrwZG0sud7c4ZYS0bhwwZZJ9mCzCHdBBslDIuCmevawUNSaORyetCV+X9g
xGxuBINrYMmN91UWafK6sDOMFb6hL8KSh7BNT7GuNG5nELN8uFJqr6tXUgRwZ8M+EWXj4PpUS4HY
MhnF6gcWlPSj8AF5b47UViCZCxoNScVzGz32WE/0yFjtYYM88GVwWcX3qD128C0Elr1n1uAHg0PO
fGzciD8op5FunMxVsOSRnwqy5aVVHwsA9GWLkQhIyHw34vAECim9HtBlc1xEE1goJubd+gPxjAYv
rDLOZt/wpQ7z/dO5IxwbQ3hUyFr1aH31hqXa/cHhQXMy1WqoyX/xiICce3Yu5AVBWb2KJVpa1eDD
aChFPa+Unju5yE9U6v2yl2QhYl9hB4/2oHpPHV7OAdpQjxlOWbl8PgbRNXBGsttCihkNHQY5Z1v2
I+De1UxCUxgcX02etrHHt8hsYrEgQNKo5aTwY0HNGFKVCTm5ckTi7pXhQdfh0N1GZM3hnwqEzcGu
R6VTvHWg9r0xpYWAY4R1/xuk4KJ42tGxRnqDh3ASCZkjM3RkhlqfciJBl242PP8a5Cvj6uMihsyp
IflqXn3lUXPUMOA85S6OuOqAbp8Zet4OmT70Hkmr4UtTBQrfteaXCYC0IwI9eMrVJgqpOYb5cUNq
RfZaNt9DYPt9Q/NekQppKmBVDB7pprHNEz28jJUuTb8c+a8pBooTnWCLA4uaKVMxJdV3/UIa1q/n
zi7rwRPUEsbLpNvUuFnxFn+GdzSviz8EhcT0A/n4Ixvpgdp6/obxYDfiAjeaR0jrkqnK5wDZmgwk
l1SiTKCZIEv6fjHDkV2SJwD1REmYjz4Sb9c/zOVrfhLg8X0RTy9PcZ6apAo81XLC0p8dyanri8oc
4ZV6Zla6jNrGo7ok1b781HY7tNLZw6dCqsQB803j1dIaEZ0s/nuuRCu7QT1xw1UpDkTOgkhR+G/j
vjl1YOlepzs/2YWAT2RmfGuIhHyGLODjdUxyv3Ymn+oLTR7ANq6+bMPklRVlNSGpJ71Q5YopiBKK
UEkLQwXz8ojrNgIqm3L2MN6nTWpA5FH29EOjy6I1UDkgpF2QL8AcHBH7X+oKKau6IR3P8l57KY0A
JEN2lD+0CIhvahafO/JPHH7TQdv7ub16b7FJi4Lk10NClreWQqHyVCo+0m4CAFqN3iUQwf0c8sis
hz2hG3+yeGL0pboRl+ZkvDh5ojo+VoOYNCL3oaLit1KFAkWln91MNz4B7emYiWGZMPrSirZMoxdO
UbeMdSBrFAOHwZibZWvvcZXirVlFE8CupANuRwbcqGnf7w2oKccU2ovrVamg+kjLBNMxX7ZHvN4o
GEhJYEBPk+vhmDX6ozUqtpJP3NqXNM0VKEKar3NJeIxulQYBJFFm/rSZ/pY2Aeniu4WrxTWSAUD4
9vcIxnlkLVFKC/Ka+5C5NxH6ACiDGjtL1X3Lvwvl+BXrXb/ggusCWk/K5K0RH6hcFuCN3QTKpknz
i9qwixx5xX/D8qpe/Tyk4uvAVooC3M60IBhuhKXAizOruVYhP+H0fL2DQm/k1JMh8NvRXj2/828A
enks6i1LOWxc2n7lg2VOAMrhP8Ll2hAuPnn8xBwizCwUw2e6LrnFSsUqhbrgFwXVMqPVdtABhJGZ
TjRB60EWqOtbkY9PuQwEnR09hJDCaWbirwSNbGJuzCvV/4gGAZXe69K2NyB6IEDa74tXyM2CfUtx
8L1bhH5Ed/UZWm88yf+u9RXwbXv75pzGgnke27oq2a8fjYLmtWq5QCmMoAta0u32iwtls0su2vRO
FJwWjWYF5C4Xm1lfmUkJzR11o9WxJiunZ73wbS2+osC3wrv5Br2zeZB2PbVMj2QKRCgp/sOHY2GL
s1zykIUUhk+ZNuI+HWow1zgQKejRAH1DjYpHBFcywEnRljkowXnwN+PC2UymQu/fW5Bry985nz3X
KZTEg42y8q2CLOvnpTGnT5rctgPPUO5LgYtM/BPBYgJsHYpgqf+horZbPHROEoIiU112HIB29Jad
4W2PfuumxZtCgrkIWQX6IMdBntyyMeeV8C27VfoJWQfPdt+o+ZKmVMKvErSo1WsUSmD5K9e92Xjj
7RfKJNXCknYPOl4SoguE1f/l1hLwcGUCxgReD8q31zaLAxqKm5YBeCRPnL5FjyMwSGolEgx1ZC7/
TT2znoognKKtng6/+YZXQT3NQ+42vsR5EWHRay8PUnhQJfpR6TABN523fXRW0HwvWh04cOaU0iNK
2lYrGBy1PLcFVmNX9orXlTjJmPoZq8+Nkvw/oIfTb8TM06ezCB44ZjwbCz95v2oPf6OhHeVtaGHe
v9VeP1M1WlNqwWMb+x2iYd4jdJdLUAOjveFMpxreFZ/iXBEBRN+hdVIEXySBcLfAPPi7j735DpwF
dDmpiwt2vpg7ZFokhYFapixy6KRdSB2HSpcjCilBPOI68hqitrB1GPYn14ybbqlVdEqNFCEoIFOL
37xXJDiJ73Ehj1KTIwGH+RJCmGkjjYhgVNKXLserexhWArgrN/3A0oWTmdnKE8MRTZnPpT3uvp0H
QPUVPnRFvvYbponoigqLLFSwW0JIbQ/7xEW591Q8pbYfjpgK/aM2ZLpPk3FwQ4HCGSg5yUWlzuXN
g68LVfcShp8Ax4KQPD6ndIQh7s/95+ifkTZQDGRVw/7eduMw/GC9ghQEp2cBw9vHGpPW7hcDG8rH
MCEJ9i6xb6Txjpc0F+70MnYnWuPkoYsTN56gGaoaB275q3t7bMTIUpOmG1jv7SwKcKNsF3M+ey8W
cCVjfRerDDMBstFDHExzTEhMETOhMZClhpFcGSCJQKUEiegHPY2ofvPcSCXIXr2hUpJ4ZMow8pSJ
BFsD7SPmHc/AbB0JvQw7ECCC8baGv9XIrDlJn/GNRMUev6mvVn8gIPPtA7f5rAdcBUeFl2L9KGzE
ssT4T0AIr+iHTr/IMVP3nJx1+PF69CokAOrcE8JYef0jXODEcrLkcPcHjGogsJ1gp8Gw+1gxe/bE
gEIqn90aMvHn3KqYuIyh7erYBQxM0sHejW39EBaH+yHKQFJZv2X+f5/hpp2pF4pxb8i3tG0M4/v+
RukBJ8rBJbC8DT2e3QhGP8/jZzO9cPDA0rHVhRJMthFDoZZas3BhgztfT74x9/k/FYkTWlqiO+b2
Ox2HJY3Y+c2o62GewC2CI+xGvvMGJUcnl2KoUEu4w+LoFMTSmKc+KvXQTwOwfzjPy3Z8iB371sSH
ObtszoWRsH+5JaoAto1Urq2WIMaI6/D1m/JKzUqVsP9ZNyjclGZ7SWU28TTtRXIOqcMZhzF42oDA
813b6VjzMu97ovmDs1RyBy4Auhd7QIYnMLndYp+Iv/Tf53obMd5z+Fwv/SOZAVBo7PCVNOiFhoMO
q6jy9JmGhaOb+NlqqhajoIkVJLgnGsuR3JyAnldzUG3QxystRz8jCjDgR+6SYARs0hyF7PzOCV3Y
LxifrZQBmqgT08MHWCslQYBMEJFO0+9Zr8xV32Jvev+RcjLM67pRyNpCm4gwQsEhEuEPJWljSq5p
ZXgy2pY93aLhfEyqfPKG7QvvjmGQmSC358frawjmvYCXeAWRlGvGTPmTNJEEIHMzBgFYAZQCR2ZY
ZFRe2UTA57mIBlDJOqVtt9oUsnxpNS8Zlc1TdUbAsSZFr6d+h7EIxYdNJjezr4FnZj/cceMLuv9l
2gLNSViwa6ldUC6MizfMdbBtSbosud1LTgJv+0uRSycPaCnqT1mNqCXMUcMLSSQMGB3Yjmmp+7tT
FydyOidusP9UEJGY/roh72Y7dtmxuHST6n96dkVT8+e9XrKW3FMZjCfjH6NDV1VXgp90Oe6IW3+f
abfm39ubv3uPDqX8KJ6gLf+mTVs4OkYhlcHfwCeVUzrsA2Ue/P2hAjFJ3KNtwzMYj1x1rYLMovIL
d207bBsKJkRC9l+t3fRTIqbrmWY+g7OFvXOQVxCnCu6hSKwvSIBqYk8ddpq0rBIrEGUYM1PcoIi6
R6LA11dR/UT0sxd+E4fuL4aowwnHOODzBve5/Mp2EN79b1zFgEuh0c60VsMLaFvpeag7Cv26EBDi
kdV3O6pmLbqVHPS30Qe0FqTjONbDCKNDPSonUWINZhJPkt1xhcr+PRVBUamoTuNYkAA7X4yg+G75
0hgetyS8OBWVAiuBH2GGrA/ZMNjGQEhboTcC4YRIF+uCU7Xn3g6FMl5HcBhVvrh7GEfDqTcQ8OWp
NzUoDKv4pwiUBm+Gz4NeVvkyxWjv7bv4ZbFns//4q/7uJDbL69W0gyq9GeB7jNGraWe5RelOP2yK
S1pvrwgt0vW72UvnoEXiUFkn0/Q0+M1/zwVvnSggiWWXjdQi+WSsX0/cRN6utSadDMZ/5yOju6jN
9SFcNWP4vwG/FW5mKwxhX9dVOg4HB/akpWLoH/REUXQDvTBnLAiup6wkvOXIhdXsi5T+Er7BLlbw
7beZO0o0PbhBD196uEU8B94sPZuX5GgFntZgUmy60ae4wDfoqji1AEcFdl60albQ48NB07+RP8c2
pk9/ka4+cxsb8B+BGBEkJJswTSNyg633+tkUKX0tKmurHL2LkqnkkizzekTFlmuZ/mcT+RnS0BSi
+0q02kaOaVz+ZPF7VnL/L+XDd4dEc3bEMHE25J2ylwYt068+xiwVzT57OwItWlQppcoovt0sVrFc
FeE4DxLeRcHofo5Tf47CD9usKylL5cNNUliIEkXHue+0+BOYoxFF0Wuf7sAqFlLLCD2jTDIvj23R
VenNcBTW3adVALdAQjZzFq9NntIX6UzEsFvkLmGoVrYaM49hTjF0FO5RwCc/iRlgr+/q6OxGMAal
Wkm5v+e44EjpShMAgrrZBBNocZErs+kx/IrXSNOOIWpcnFLdIjb0rH2j3D8AOmIbUi+k+9/UpPuu
f7rfXDunmTuSfrWrFOdcbh9QJfipZwaNAX0KRp5WJEmQbHJiNvVN1nH04GCBPnZYTfseTiaUhQK5
zOKx0CsIk2wZyq9YLhu945moLmnM8pDQ621wlDLQNW4z1zPAwDo7IzMK1C0BXxvVXhC+aYLE+lDf
kQPZMV0cW/k8ZfXHUK3wYKDPfOcNih5mrVUTUqloe9csZDmhMuX4mrWbG61eMyQsw0CCjNbo3jLt
9TxOxHkB5MDYaLTg6QduUeappLSWO1+9NL6qaved2ev0A8JtHhh7a92riBKoam6l82I3qm3Fd5lD
iafClf8LSq8uafoILUoHMrps5fRaMTLlbBlCKsdkIejpwXNmo7TosS7eTZgV6T9s6eUyut0L1CYf
iwJBnvAh2Biv45/2ucr47wTW1ip6WZ3tUSqYLHmNplCSkoQy9lAOz7yknlcwgfpnFi/56otGuMS4
HwOO1VBw+Z6HPzYlQPRe0lZptuYIZ2kZnr8N7JsHGiKRBucFqzn4vgVNjURKhxhHMF2Qg+tp85p8
uIbAnr4wHuIxVaMbUXDccO00zpZ3f7wegwTFtMfYSInEsH8LTKO06YFt2xfrCEs8RpIYyOGaoh6z
0H1vezj/Kd5YHDkvW43MXamsFLOc7/zVivIzuOxtI28ahO1fBBk11XujOCsriO4p6ZT+k99WDsaQ
BDWohuA1e5weKDCXuFjG5JXdugyJGDu4Vn6WbQwh860e7mVuizqJyTXKOYrDFyxLMHnGlcH1QJ7u
Q+I0GhGbExwDRzfBMSUrvA6vEyVb3Ytmd4nvR0iFHBVQG+MXsmBlj0wq717s8dYi/qLshoqXKwxM
JC5Yu6r2wqRKY+tWMTLXVcNEPV3rl/b3T/rJBVKhVpnZX+GglkHQB7APcUJzzpnbDvfrmZAK2KuM
Ox3Wzn19E4XxBbUmML498lZWTd0djiK8vdp5ZeU66sekZWZnu2QDqD3pSV8HgVRwptUG+87xq/IP
iF1Z3SY078lPckttvCGCi1X3ynRekb/UWtPQRKefk5XZQ9r+QZlU29d55+2IPULrZnth1teA0BGX
2gfRQHj8aRpamZMlSFOJ3WB76ez91w8s20XH7JxKLRnU9JBPFqgd+2iVjX+ndIDlxPg7EjsGiVhL
8UBsawAry4n35Zt8DK4zUbjtArpmH9WhquFSirOBs4iboDixZaUo65dTDw9Lw7clSSGtqSDUPeEF
mPySOdH5zXkQ03gq5aYellHemZzM9JVExdmCJ/z6HaYzCcPGcZLBLY26I2B/wq6VDgOT9yfLPJMl
t7UTDcvaAKqfz6a/veYc1sDPsO4O0IEMJgcde+ryR9c0g66/B/GZ7fgVhdZdodT6fpUephVVAgWC
1BoIS0OLxmbuwV5/6zRfiydkeyzC0RAQkSISvThGKMFPmwk8yKmZE/Ros1sGNbClH2bAUlGjeOBz
r96ND+sybi1J3Wi6GqZKYTtG/fzNJXs6xTdjo4hCRQYspa9yeHbbKCxxfTV+VoyqOubgm35HMfSt
mRCTsLGNY/+Vm655Wvwzznkl8sKj8KqYf+6iz7fZ/zA0zlPwgRNs+c4DQghhSt9hZ3REwGGgLHQT
1wJTCZED0WCS3edOj7V+miU/wG2bC/7KjSt8nEBFhbPB0XAzEuhLYCYQwGzPro/mdUGhCj0XVtHe
VUNHi753NKYeq/5MyynejwGBa/Cx4kWQCuKZscP3ydB34PQP2F09LSKgDyMRio2Y1s/b+INN/cSE
nkrcFmakr/fks/mmaIj32NC0izOesbeasUSEgZ/az3ZKRtpuhTEkHg3st1SHyG/pbSt9rE35pnti
LkUjkj1HhydjfsOLEJacRPcuOp9TQBM4BQL5xnmS4upJn8QZEXjroQK98gp1NxdHpwLRWw15x8s7
Ss4o1ktiAqdmAB3IiKef84YrYK+3m4vfw8NhtThJhoiScY/F1XfRM6k1mqJKNNf8Tykb5rQhF0J3
Fqn7hk0fZ25IzW4EHD7KbuNnFgvFboiU/ZfIdfNoALq+fw4+znC6ofCceJgD8X6my+VELM0D+MpB
4PVLpvY4yZw3JEymFZemgDE+gTa3xTRxFIpmSM26EORf9z7umUbucFOFlzCOLoplykA8q2YQjz5h
X9K8I+hXuhHbmQ8hPbt+NWNNTl0Rao1obXR0Tq1Q2Y6EKY8WbzWvVw4F+ck25S6QYMgicO/wSn9+
660FS/TD/h/bI1UYbsB2ecksogaNfy3HUXZQYf1Nv19KmHdZdEAXjJ1so2pDtgm3xrD3iSPW+CWF
IDQuGt1h5/r+ecUNoTb2Pf6d6VemiGerXTho1slWlXLom2RrSKgQrohtkdHbm9QFTHwpbtUUgVPg
ZwA9LzbWx8Ov6prmELINwCIV8o08FjbX8928pxtZ4fdoJmocz7Hju30NZFTOneXZgMsgHCbEn9rD
3yfHOby/dg0GM6yPFpYZoTYqn+7o/rNx8VpyK9oLcwL7uXutdD2MJTCgs8toJ1ywy6pTycKcheeY
IkFA3WX1w+UVd/TNL674ZnOwUQKYwVg9S0P0XAslswK37P0xiBaD/AD3LmqBCWfjwMeeC+PXCAkx
PH2Qs0rfSTm6uzpbGvLcrgEJxLXMLzpKGNv8E8pZy0UyZ3aIPp/oHcymxp0HsIYe/i9dvCgVzs4e
FidakndWhqpeA5LdGsyPmaLl3WxpAXLykB4VoLz/uXtz2z/yPsE9q1Hr2q7xWfQzKigBR+JNNol1
CQoivOQLAX6okfFIUM3kD//XZ9GXmCWRENRTjy9ZFl7DHVKK8hv9AylVFo0zsEDFuUltBTn1g0sd
jmSg25OEffkiPPqWFWFgMO/lHjeGQFh+RRblbVUD6eJtcfxUkfGPyQilADWVEMpT+LM7YSWQ7+1s
yMjphUFkeARuAl34UJKU+eTOcaih7mtshnH/AfFh4pjJ27/YH0KexP1P8CX8wprNmD4JYm4EckB0
J4Ne/E5XXD+ZTQPnhaSaJPZjIn4wHiC1rtYbRWxcSoSNcM3Aaq3f3Hhz20VOsBi9+i2fc+8xxdkM
ELa2lG7Vzt+47H3lgf3UYce/pLZZhsjTJXcfaxx2zAwz563noTdE2Lf6ZeqATVfgbj6/9ddE5a99
msBVyvmxB0mEkWCtEGCveZ3sSZiXevZFEgiFW3lpw8XnIzWuk0ymyaVBqpcaSpIhqfbvxPbz7qZo
icHvGigsWPMj/qVasJRsx55XC42q8ef2CUR5YRRDbg29LdwG9BRy8odCm7CNiogLL64ZAfEV/xcS
ZnBesa/rAZLN1mz5y3QJXa5Jw+KCt4Lhj72PgqlBO6RcYLPHkuo+/r/zqceIAZumZ/qMfL9SxHDE
tg4sd0b/+Njzq1R5H0WOoKrAHNrmXiakHOn7MU04PIHalYiu0mLQ/nO+GOE/rOUtwkqzcdeKzHFK
eKfS7M/a4Txae3fhnuH68BtZHwxOSD39CnZAwCB/eHd6+Uj67BVCuxNUyuednTaQ1gZsJ1Dxiy5y
B6zbyixrhz1UVeZ3RiPAibHhVaM/4Q/ciqxjhoRvJP62m6mbZqAWTuU2AkyFAbWACd04wUUhVdG1
kh+z9Iv9TbTizO+nzNDgw2CmdaOU/0mnA8pTV/VaXvdP9WKXa785q8/OpWyn2jiTMjPoB2WOiX+d
Z7i+nS9nCj/9xbLobfx6jhi6ahf5j0jEReIcZENCiWuGf0nDFX7J+zEf6exzb2xssWeiemykFY2D
rP1FclvU+jjYC34LP6VBfIhy7GPDGdAPSXJDRxmGvmSnWgxOXH0x/UTG5UznaIIrcN95vJn44i5g
Hd16evUUon/uUvKujIbcR4YuFytEbwUmLwZqYcAelS+tpftCFeI+nMN6rOHjwSMY9W9iGXM2Z77u
BxEjbT6vqPu3sq6WW2pq6aQoLHZfP7JXWQvBucsKs7T9afCL1iugmHuuHldZCmozWL6OhglZhDYp
GvYymBQ5GW2KlRUtzQESypa/3wPOMudkNltGoULIAbCfm8RhfpbYvi2wcus5jmVQ+ETHYmK783+N
VjsMchtBaBeaYEF9APtuujdUN0PRUadWV/RT8t8GLHkExTlT7o3fApR3GURjgGCDDILjS4weGBbh
Rtb7aJSUvvJgZrLa/KXcgW8l3md+8cyRQVkDjq/kKXn9nKwvE4pAHlPnlfGrjs4BeJ2/3ia6wxCl
s446Xg8AVQeELt5uHL8RWJv3QFOU+/v4jVEVuXgfiyc4ZAVGfrUt/YvhVzYUtMhkZylNrdOECg6n
jOGkqwBcsk+1i1A8fFRsmim4krWZY8znSUJSaI/RQAoInMiHs0Gpw1cjUnoD/jVmgsH8NOyiSQJy
9u05uiJQjz+TpWESuFYUiSEHS+IkUoko85o5w4o1ZqLIR6RtfD130AtbKEzj4yDnkOh+OIr37abs
ykwqiLXGv7QN6GoRE7Z9FinREYxAIs61NU/TbnJf65uw3cBKMFY2RhWYMVxd4pJ1aQ6jP78DBqxe
lt1P1iTOV6ifWZ99DHJ6PRF007zfuNAipllzVWwyMCPWMKTh12/wFrpCWsKIRz4CvVW5Y0fs/M0F
87pXhA6Qnl2VDMR+r8aH0xTIEFy0JnV1WOoHTyVnbobuh5TbI/KJxXxjfVhGTjifXK2UwK/Jm8qp
2nEn7n1/+pgSlidu5zc7W1A7N0pgM992QolQqlcHeafRWkUyzoWAbQLF/SDJpUgjW64kSzO1WIbp
fn7jxSEfluaf+8+KvtzH9uDqZ2n0QmubvO3Pm/GBmE3gjKTl3T3tGzlG4fKFe2xYALZIQxOWpntL
4F8ZaLmq6BmmG/yzi5H0SyqzhI7vVbLH10wIpSR71sbzIx3RyCzXcOxCaKKWMiIQ+Q8l5LhwaWdo
Asp1DiVaRMZV6C97hbAAvvHyuN2HMisiPK7ty7va8If6d83k5Qbpa/ZeN0cLM1fAvqtyvftWpE5l
kA4nPAi/6v7TpWs64AiPxH+mvl1BG1zPYj6eqQL3b6FSvTfhNVKb7WxCW4MSdT6FcBmgk+bd9aQG
ElZjw4kUYTI0E5lXAGdOMFwlEZ7wru9KZOlWwtcYmKPawEZOXjG/n7CEYvXTjf/+49d7rHaKosId
nPMrrq/KHLwzE8FsyRjsKDNyp0xvae2CirBk5ZSjzdnQ2zhmjuJgKBiwa0kPFKf+cTPcTt9/t08W
OXve+elBHzauEqHe7nD6hl23FIDU/QomGSi5kTFBmvYFRA0PbAsJAlGqgOW/A3prFm7RZJPxxCfp
5VK7PF/3MYme+SwcTO1urTlsSOViabEo9jmGMXW5RmH1uKSsasgkYmT05gPq/23OFu3W5k2Nf/nb
TR81AAnB5leiFPu+EL/ikBK5AENFnX//QqJysFndjVKAWAVRppnxwvB9xcz0djIkjUNK+DFO9beb
xJWwKzySVrM2Gl9SsgaUOOM2D8CyqOQeDUy7YpQyx3u+U4macKMEuOTkGJyzYzSVqpyVzsFRoMAV
xTXMFcYj3ipXFPgitHb2ZcfGWjcZKAmnr5gp5s/31MW/UaCIpulcBkLw7eq0vx7lHlET35IdwHGY
WGVHMHkv6eqiA4+z/tMMuYE/P3NIVIjhitbCeUdy4L+eJZdJhBRG+qutuJk+T5OK3S7X7QG5tSbC
PKghdwGjFHRsW+6ntJOuM9vZBCr25jCPRZzOoOXV6AN+jlqkTJfU1gD+ZEvGp3EhcnlrBw3gemBV
PfrVmuzrZIdip41npaZLSoevaKNaGT4mUDEE0w8Tw4xaA32fEXCScKnX9FcaWbJc/WGCIOO4IPjC
XZskmSGIsiReHfWSvHAJyVidB7lfikyhA/wla/nm2QcuD5Bz0OERPQ8h4nPPQ/F4ueQwUNBDe/jj
MhsQtGUHSoIjMiNkOkhk2LORyMtPcBw4SPRtJyA6ErnbtcBsiJ6AxYejXElCE/dLQ+E8rNJmBFt4
mwPicLj4SrKpbqSZjMG1kQiRN5zag1S4eT3ueag5t24aNkR5RShNlxja0wEz4tnAUsB4hjktUNKU
RWhxYFYASq15s739heYpqoFQjapaY3aHbGqUj7jqhGyDr8ayXSrARAxvBmkXYvNoibMHeDukCc+I
vQf6nhCSij6HvbFLZU6PD0MrzPJtxCKeC4iySkI4aQVFJl+cYAtRj1tTLLizIm7TZEg23cr3QHzm
5Zjla9Hx/kJ/MlDl5SRaie6U8TK+EzXfFLJo8pSaLFzMzG4/6DdxZyuOdo9Fe151TMayL1mNUoZS
YxLSgEg+k34oRwlcgeCVEGDO9FHoVSfgKLXY6Pd0qv66c40qtTvNb0/YxWCwdxqheodn2UY+iAp7
dsn9kd4aPfViUSpt3RwZ5ABGqaNCZ6cJMTo/PS1ZcmXGY7Ru8LwxU6/vCVmfhtoZmxu7nsVYl7EC
gGl84WkTsgrR377er/XvZtnFryZJxn2ANnvzBuVJL9SP2xvBtLVcIeTFLlWqZ2mLvlVyYNLGJMxb
7G6kHelPdhqqqqlLFaZq8oEuG3GR/I6Q1zk7DKQA+qV4T0DhYW4uCFwYhg8JKVSkT8EMuyWr3tFl
1uYi+I8kfW599LEDhjlpjfLF7mrr273QUCYRBDEsdeZg/W6XFRkzj0t/8Gd3qFRQ1crVT5WaUwj9
B5btkQedKJ/MKMLKnGJ79+7HmCsGU/uY0BsT5OaD+GBx/VwfsaU96x68eIpHg73AsmbHAilOZXN7
kru0/b7d6qIFWjHXo79Re1LOhb2KJO/Nhd0pIJ0tx8jT8A1NWP+KGPA7lJb0McLTAS71RIPIS/Nc
3nAIPMCFTVSnmrFm8zIYwjdyOfE/B5fOdGn4u88YX7IP90wfznkjnPfUf8eQGsjkDG9euc5lrH/m
Orun0jxABJf5rDzJIz31+vl3H2t2pMvqov6NlpnFc+ouukd3OqxodSqUrzAIO9cTKyMdEbirdFn+
wcO4cHk2LL6NM0Q27bVzy0KMjR8NlN8TVgCow7A8oQFoqQrLeuZGogCfGzlAvjlZtDJK2PozRtep
9Bq2F374TZM4O9w28LZB/VuUv6814pyGBq6ePqlmL7y4Xbb7SWLdHF04grKPraNCoKX7FZnn09zO
nhGdScyMP5T4EbGC3RqUN7ezeFQmsEFdjVd0db3mSjYW/oGLtlF+GoBifYv3wLJ8qPbdGCGrADBU
PAgbjPY49qmHpUmMITSF4MsVY4FMzEaZLF4uWz4+rm4SGHYN4IKVp2CmUuSHPTJBbT3YK4op+Ykl
X6VnEDawYNh9UVZ3/KQxlh+KW2yE8cToX0FCPiAX8K2Q58OlCnGeKZ7KFBqk09Ze08xUqbRt1j/o
WOjzKv2jBsHMaxR5hsGfgYZCBPIwuDJOqRGFtbj/mk3Bf+790njSxFioYyWC3byqjdLLieBUDoFv
WDPGzU7pDajgAYvF5UWSv8qhnveEH6ro94af0csXSX3kv50z9/CzbyGRDplE8Ul145IRG7Z+9HYP
BMsNOvmrkU9z9+FCQkELI5JLE4igMNXDRiQF5IBNWK4qud0jpFLAB6KMIYUthQ065PLOOFIYfSSt
fON/SDz9ih/WbuOrXdyy/TMb4WjgXSG3gZrSwRKYReKFh7Bl/Lj6DDs/8MPh20qIwCymiheX4xW/
klROAYw4qyR6Wg0jeZmMCa2Hn3rHRhAqo5SrGdWMgjvv7KpzbKQVPRMMRZozleiWn1SCzpA63BfL
672t5o0MBMIQ0OmpPduP6irvZNyB1e9wB3OldwXjPAgHL6/X775O2aeFSVCwEMXFeStYIWwiZgyc
fVXR3ae6vU5utmZ0hVjLPeonsNUpxsYjRY5L6L+LA9/OTd4pCU1OZ8eoIEAMAXaiRS5tUgSBiitT
OlTUHZ/jqPZJEqIARTaKv5vseg06BeLXKPpzqMr5kOGc5yoxEGI4gGqtsWFGvedRYreGaA2C782v
Wk6Z9/7uqngaim5FtfpO7WLy5B4Baxg/S/wZAxSfoBkoZKB0eHRHoE2rSTOvUCzjfNYIpYlc4m+q
S0Ce1en9C0dIScRM7Yj2spnbLQxN8PDNm++74OoNJfqRB5O14IYANRBnVd7NALOgkkPTd5MDYsTN
/neZ8w3kNUf+Uv+gNHW5alQr4pYPzfRl904CaHj23t7PKZMqtQQ6jDUt5hLhiTl8PRLwssi9nwxY
Bx6Zd++mpGeBjgxuyWtK2HOZSAtpu+Zg36Au11eyOjObGOhyj0gy5gaT+6N46kVzmOQubqIyHF/l
k9i+A78oFoDk5KNYaIt4SPlBhEhy1vDHxgJaKvliKxg7TiBIMXGxpcMCXuB9ZvsJC8DN55YCfrlZ
r3UPB1wUx395t1bPLtdF2K7vHrjwsz6r1j+0AbJX4dpwVC92LvWgI8GGby6tXDuo9gsA1LwEnXJO
ijhd62u/ziBriQhUaAAV/7BbNxYaTNpJd96bP/vMH09pykuy4//42ciDQWSsQ6KVqV3P4VB4k7l+
a8Nsb/OMWAeKRblX5R4N6osaH5iO83/5CBMwOKCrtgo6nuxbvZhUTlsOWHjAq+K6aOFXSWq25xkY
+l96C/aG8+7IW5rLch8MtU3tcgIGHASbp7cVDORqg7qatx9PvFrathSfSzXDPzVCJnGWDMODas6j
aGX5ov1L0EpwkCknlRaTQlnfQek+Jyt0s50tqEo6doi3BlRbaRPKIWUXNBlxUOzEHoBw4TwegkqZ
Ubg4fkx30OdHSpaDyIjJr0PBoAZVhyc+Yo2/wuFnm2MlXpzvHGEQc+nkD1R8nSgWv9f7OWHUN54W
/D895LTp+/uUBvrCf+ybhsqyP1Xn9I+SAClZR3cBBs3/EfuVO5uBz8Xi35oBgcWmQVEXhf5njbbY
e2HOF3aGJq+XCKknkQ1bH/UMqeNP9PeVAPhAztjV6icsKMkt3zF4s8w6DCILdjlVjCG63i5Llq+u
meFV9CcF0SkW40Hffe9WlbD/9iSuDGs7oKs4qUK6ZxXcZVM1gzNPRaVl786YqmxUZacwYCazMVmW
nVy5wTSnndSYXJ7x/Xw6R2KZp1IVpX18oixenBQbk6FftUPK5nBogiglwQ3FYJKa+SSXn2ZAHamI
KDatvQ069MGFC1GIgSrTQLGEMKKVLAdHgKijqJM9U02HWw1my3CwLxODkDly72evs24gfC5zHl9G
6y+57QqzV/0aHC5jp5ETtF0hWROTjnzrMgCHLQ7cN7xpjx2F0pPhWLTDgGdsQKBZFvQKWWmKyBLc
YpaTcfvYshU/rOgC0pYRm1di54j9ukbrQSSirrH2lhjmpS6XXrvg2IaQaKrjr/bN+Qrb2WRk+iST
HTmYhi5We0zz4evhP6iEhPhv9GRFrqRmszozx4CLayUX/qDT5r23zmNMQEC3CD5pnJP2IoXMeCnH
Tpad0NAezjS5tJKLYjv8PohptF+aM1C6OOqsXq2JBleLJ8lHzHaSqq1AlQhELEnNzQuMchHFmI4R
37cdzeOOqD6aHJwkhIlVZchPOA9+3lShoha9cIoUG4uGr1EK1ep38/xKh+VBRM/JgcFfiSMxWRlI
CoBdrqdLuGlq+yE5Ps9jM1pmWsaMBuQtWYKd5YLxm6VIIfki6FoQkjreVaG5zjVIwnZixDZD862W
3Acg0hC1qVHhaDKZCY8DmRb59dd6bUwrMvSmwlaixjlRuxWV12Quw1FfgsMAH5uX5F05Vdo7npMS
eS/zzUjGhxACJstWxJsOZoIlk+BEZaZN/6bPyp5bLD5ZUKi7A/BvQjxnMTiumuC7Vthzyon3SMAR
B+2vq3IyVKmC6AL6iQIzX1jfiGNGYmT9X0y2Ji2nMKrt/d7dWbRiBCwo/NbT3KEdWwZiWjAEfX7C
xJ+Zd5KvvIeDa58fNtcBGGv8cwSiEhgsN4tKMrUmYS4gnn+lPl/xxfrGzOne7cgT1Q968JlH7XNo
cP/e7ulvJ2hlg3bInpdv934dtMS4ig8sd8mNn/3+YD7gIXsbXbfSbu83mO1CmQL621RhSi9zUX+0
LUyxU1m6GmdY6hnDpHI+dJjDrr50OKonsUGVl0ne1cVnon6UQuVlHNaMJsvIOr0RtA/UEtFmxBhJ
vdCmW/ktfl6rAANN/0Kz1dscryJEdkQPDpy1F1PceiO+wZPJGHzec7ibuek9Zi20bJZJ/NH1q1Ps
ZywSJ9U5PYi/Jxc43eL/Z1CFbXNmgzWaLhJHx1z2gPnRNnzVkrMNEy8CI6qUPQn4k5bb2GvIOzpN
Ax/cDRC+vPWAimoLA4WwZuwWtjrMrz2gTaGiDDTty2QAMMnhB9CgJvbEV95wLiwgbpv4kCYfhFdg
BMBvTsGbI8gEPzRPrZ9KW487wFyl+nCnQZxbHflHUPk/7qbHx7LyeOhj6QvnWOEMqUdRCx7nI3/m
sTU4ph9U5+iCFp4XIvn0Leu1tGa2A+/UhWyJg2JqfGo9e8M3M7OGtG3rvOZfZbau0MDNGogh/xHC
X4hFHTu2BStMPMezO7jpLRjV/ld+d5GSOSxxgDHd+UIltVRihzQHUagf1vrgTMWOu+EoksqZEQVk
HBAGtPTt/xtTRz4HobabbS6iOgcgrXCGhu7Zjs1MzkZnC7IWCPUGR7O59Q5FAtqj4pqnfVrj6Agy
HQ9mj8MNuw1PuXvTj3b/FHst5csyCq8RUES35xw2KP+wg6i9pf2fX7gwFLpMF5u+G0vFKv1nnzu2
RP/IYOetqmRLmrUODrUfl+zCPUJkYzL6nCS1udcw9FwTwTTI8G0ln+Cvmg7htOGva3Yick/tkPWU
Ys9Jw4PwVV44tfAQ8JkA7HFVwUcUiNDc7DI3jgDB36USvn7KJSx1vZ1jLGFXXodnPhDyb4ASzy4f
3a73yzCxNWY92bBpNS5Z4ZQHg4A7a1XUkqkLEseSwt/uW9Y1UPpU2s4/8tHjni7qDClYvTvXL8pw
Vb5ya50CIbxXANl4qaOI/kQjNUiwFNlPGhsY1zG9/nzV3soqCShiY167IYWVOQq/JVExUGPuZjMp
k6DjDbgv2Y7lNVj6rkTWzt8Eu8X+q715cnHvpbh7UpQxmaUZFv1xoEttht+1XWgJqBuoIxUuTtdM
gcM6ZHHPQCChXUXoE7/OCLwOd2n0jWsfxm9opUCUlkbevupmbULUSvAUI2cRzUjQ9aV1cIl280zm
KWDu/xi5/B67p1WByEXlrnvI7U2YxGj6jpPFr5c5IplxfcN+sinmVDy9gZCdyngrjZHsCKI/PBt+
1f88UvxsCjcHrnSMEzsTQ0ujixrcVvum+c98wI85J6K20NLsEXVjpKH4ca9mr0d35YA+klG/pKmU
7SQrPOpp+BLIbjCX7/1NB3AQMI/XRyq5PVdjkHgxv9IJ0KSEMeteiHz5I7qK1BjjUkN7RPxQC3Ac
wfs8qMOYlufa1GGzqr0m5TlrGf8YTsoVIwywD4CWjYDNdFWnG8jEchsLiipmD9BGDiO5fwEbl6UL
q0zoo77cbZtBefYU8cKx68IPoKCf4U+8Q1vN1PYM/y/gvrMtaOFHlpIagOBrd8ECOxuvyIJMSCON
zaTXaEnsQbkigO3Kc5WXM9hgDsjQKLOo+QytDTD1KBnuHxSYS/lz0dmoyKFVbEGfBqn2kCLJdM3g
uhfQdbN+3oGUKWaMa8Ly5GlLEFGoI0wIGY2pfL6kTf4RaECCn2ubkC62A8t2ftoSiWpCOzKTDazn
+TvNI9QNlFilzV0SKc7jIijJt10jjQnntLRrwX09JgEFXHow+8JnJhtrpLsTEPXMEN3TdvzOGHGb
80shkLwfn3D76O/HFPbfpnHaaW+Mw/gX8pgNY8vvcHuDTbG9e5kuIauUedbetPxeTIWEttCdEBnz
AW+UyiFYEqqS20GSJW02uiQrvt2XniDqZ9Yyqo+KBTwHPc9OVZR4tUYk7uaEJFWQ6VKnmWyVVeS5
eb1HhtcIPFlOsKtzCAlt6fTBgOzEvRNU/gkR1D3jOJtnd7pe18jD8wqwGDHoe61ksKFg8YLRmxLp
2YbFUhEXAVWos/9wcR1XELSjDYWT6FSrQzLHkTa/TZXqqBCQ11i62kkN9ILqnZEHIBCkqMAsgaM7
Lm7Icf76XxXSvnkOfyVOY6B1fP8Wrm3q/KVh1ap7m9cAmTX+uYAcwK2EcgTy3SBwoYyiU/2dMlv+
9+3/fYG++a6KYFRLrv0UlSOd2lRWcfdzFpV0YM3faFjyI0hmG5aRVUqsus4EzKBf83NiHlDIR9Cz
OdnUc1H4E+aPxNFQQCiv7DhwCGuy5RngyxHZdqCxJlOVtwBzeXYk4IMhMGUW02ZtZSeKGibV8P1w
zH2x3uaAuXaRu49uQMljrmVp3iAUTghpninLDIqp73q6jkx2TY+tKoIlpZ+9ihGYlbYKvVpQmPf8
90PBhZCbdG5JWOSMiqFIsjz97RG1pi2AbmWpSaDQNGQ3ewI0yyFrmQDcPj9pTn5ybU3ICvTj9ErK
+6oC6KYmAGAPSOxWwR3wnC4dlQ/T6pYxfU25THKmFS84nTnwHpA2e5QHW7hM3yB33VsJvcmGLtJW
ZDGHefjUGuCElAhoUrmxCuawPcKfwujMKQbZ3/FcbYYwE8Aa+4wG9Kp2U2REozfCHw6KLZDUZoQf
rmh+6wGYRLccr0k+074j7cfoKuo53XTodRDDBBk67HL4GenHkKVEigA9l4ETTfBEV0GY3mslwbCM
jTJB7BU7TGioa7Tp77YuZuG5g5jPMDmAqjwEBa0uvNIuc+ltXSFkE1v1MMvldhNnXBtmYqadMrxD
W2rpY9wvOtCtH2KcJP7VLG2CNk8olZB2UAqdLJSRiA8TcrF02ynMJlkOG3DGH0Ic/CFnTPCqpUw+
vPdtUpfUV1rA2Jvodorz1WvPpfnbxJHt/2G9AZiYeZNSDtkhe+AcEecF2cBlFV+n0KwkIKlp/+5I
t0s0o5h85l8tKtvPGvC8NiS+G4gZ0A2RkAoh9bSVbnxVlqlOJZWFhtZjFQ+fzeR5He2oP+xQFazN
49S3q0Fzo+gioZ05wO8I49AqLQRdDZ7LOnlkHPHcqI0huyAB3rURthtEW/cYOTtHBYa7SpZZmZHr
q81Bprt5BZbEkq8ndAROy4AejR3w7OB7vptpUwbKM9GZRuPS+An6tF6AyxA/9I7IUk3mpkvt9nVF
d0OzAut5yfSLfES7XpD4lOLGAB1NrpcscOqvzBo8HcfB+iVGoRy6qBy8DtfQYzQWNqNUxF3MheGI
/XZKsKIuiXvjoqC3m1VHtKZ0qr6/JmkKqW6brcplGvKRrH9e/sDvoH/eeSCevB3iUoqjSkf2jRUw
sxnfjxEYuP6b+y+i0PxZIWsWjNo4ALdSUc1T9oPrP6L6cGQcZ5jHPZiSOovcszP59x8itkjKiKn/
gGb4h4faKv2B5ssbYGNBAO6GACBhp8j+kpgPGtdKQT7Iq/V2RQ7n+b7cXOswfxbS+0+hEMn0iYQN
4ONRkGQaWjbtuXhQI0cfDx9L9hqskBK3Cubq4ZIGN0412rbt1YskrYSgAwcJJSJMKlOCb3S/Mtqz
bJ4++ir59kMm1/QH9s+CDLrZP+SCbMC6bMaJDIu602fpOZh2hHo1NcNAscsahL+e+1fM0zIBbgRT
y7Bxs52t9jRVPgT8tOy3BW3HIgcdI/45lwbMApCn6CyoDfXUdhiuWV6tXK4ULOLtjOAyZvB5bu7y
/abhFEFrQFc54zIiILpJST6NtG3WjHKgz3Jqx0qbZx6D2/CZ6zQWKQ95mPvuVt/yvlkXs5JeO+8V
AIq0MasdXsErDU1HyQ+aNiVfiGLq586PZ/LGJl1voINfbBk5bHZp0PLcgOxs5CVoDJqtvWYMFLPx
cCmSGe7HEroAWH1X5uzKaN2TUKmZ11wep1p60bQts7AUlfc6qKqwXii4nSfq1r7CBL0lPqE2lBRE
kqNL4LvNdHM+UVe5YOn7+ofKQClrZLM2oYidicKG3nvzxtsrTeY1Q7YEutMHTARFYcBNO2JwlYhf
+EteE4D6M4Al8/80MUQf0Y6NH1aKDXHJFhsof36Ei559epMef38bejSxDw4py8kT0htQkzgtzPLB
4uoolxudBtaVa+7lzBTwA/ukBh6/hP/WpanOO+nT0qcjSkUR5DChRS9IrExbB76QbGUZB23Al18R
mjDPSJPWum2CxRU61OQGrFf40FCWOwKkthy1r1CGgIhYNyHLRruaHhBPgCUk6eZbCEMgej42+DFJ
C2NcJ3Ryr0nox/1METx34FKGbN7zXcBMw4/+R/uDMyDM9RjUay0g9iY9HqAxQWiLpc4ewjPejcwr
JK42ADtdaNV45gl9CAZC7eRVPku9w1N+9nfhUKZpARNlTBNJH9iAVjodysnapSWj5fybbmmZGHvc
2nQ5EusAbM/Sf1Bq2QOKEgLRG4k3jyOhHb7sfVedONHZMsiLy49tp1keTSpDEpaQuZunqtyO7Mrx
CtZmqRkfYsRmaSS2PqjA9WPE+tz1H4hB9TvqNQ1y798zLXY3F54PxD8zHRBHPJ9mtv3Hxar8yAy7
v/KJyE+HtMg/iZN0yJnldthx0j6EVqUK3h9ro56RHjmuX+C1Secv//vSbK97OwfE3K8FGuvk8e+i
IrGYGzoBT+pjG3xZg0kOUxm8HpPABzugP7wWXoqqAyXQWwtgzcBE4ZIGJo94Wsihh0yTsYhq3JR8
rEKMA58z4ZHfTQFdLr3DDwtETu7aBwRNME7mPzfpWZ5NUX6qhuIztW6koDWE3yVZgftrkM3EvQ09
lmlDUi9U5QIK72bBkpyJzdDTEuQbYiexBgvfmC4xAberGQtOQsWCIykuEUGncFRN89lxxfB1ppjc
iUmnQc7X4jwZN9jVfEVkxkJKSJTEjC65ChCtXg7PlK7w9912IqIVvMtxQQ6MFjTKmP7ofWFDN90N
54iB1p32YWCLQw4PVVSC3QsHbSncEXonkD7TLlDMWSx472+kRBKzYwxmLr+1okqoVJG7TyVlMpIe
48OP26+wG5RwBBVsik+/clQ31JF7Z4mniiPn2+MpSVsEGDtwJmbZDGq4UWHBqPBhQifzGbjw0KQP
Ht2Q6jOQ/zY+MokcioL4OexlwVo+TC9bMjbamNCZh5haf06Br5RpIWIAq5LwA/FK2nnNuVOCXIaB
vKoLsJbRwtJ/V/8F3pEUuzclXrq5kGhRP1XGcuvFyb2dkSAFpZbtK6r3HrIb6kksRp88GGMtsoHO
1/vpb/prx3CcNfiUXR8cuNVFDFXk1UpdttvNrdi8bG3nuJM4YUtbwtimZlAyWS2z47jMGhzjuhl6
6zTvLyUYRymhcOjI8VE39MTHmQCBAwvMfn11ebJVZ1sthsf+PSmAfD/4TumaUf1XJ2vXoPoH31mn
YmzAGseOlQmj2rizzj7cYZFgikCpf+d3MvuRKt6BL0gsAFPVRDowSpSa1/GGXzvt9seK5bmfdZbZ
T8oCP2DdIotKSaUe7Qjtfj0wRon1Gbmyi8L7vk6EmeS+ae/h/0gxMYf3XR/cqBPFEGmCdV3AE6Vv
gvz/jm52+ORE9YDxdHR83YZlR7ps5ejspiPMRCKRoii2K1jYgj42JpECqzTyYF1GDWOJ/QC/+MkZ
eP0m+/ScBVeefexKOEHKDcHuPMwsaeOEdu5GEMSOBpPYsSuMB+6uK1Zo5WA9KLkXmnajpIWX9j+i
rRDcocjapA9rbAR8prwBuAq0nWoBfDj8bfPcxja9ZimFivy7vulolo7NDw6rK2Rp/feAM4ca2Nqv
OmmWrrbhjCXS2MJNxv0+bCnX4gzb9O+Xhfm6ftV2blJ7WnsECDGUonEs9stBhnmJut7Y6eoaqxw2
06S6q43plgdffWBCrcQGn5H/XYPU31VrcDgRR+f6jwv/KlYreDM6eroKazpPcuwPHjfLA896d9PP
6F3zKhjJ+XtE9nt+P2CZgHE9kuVCM4ip4w6/lb3l7nnhLrcO0R0C6vKKoq/KKNiBOsqvQUnMFZNx
BCvub2szDCZfmgq1laDkyLUruDAsEGZZx4hAxS6Ns07k7nj1Bm2TeEeRSfnwsScm4Uz0JWffcmuk
DjgqxJ72AlhwX4LJJqj+5w4m6qbzt9lGZChFP5sd18gYfMlyDIgjlL/mLr3lt2UF6c1HB13vmO/f
ZvfeHffjh2aV4aNRfThJOBwNfhj7dJjEyfGltZde3vrPNWgnulwyyYPpviBswYpH5sZotTjL+NJA
n4ifbpE2+4a6nLZEiu54LZghmijnMjbE0lls04fnH2FmfXlSHwBruoPjjOkx0G2e3Up+rolhRT5O
/b1RXds9qPcdmYUf8QZjk9tPRBwECoHnhuK9UYcLMypjyy/KYXJJTho8FoRyhgXeI9bMx3ChlXDT
g30QLLF87vi1LoGrlShPj4Hs8FNLgKLyyZp4yzoPkKimPqj2coygK7FM6CuDKaE1N2xDy99K2Yz7
KeSdnDYUemhPJR3gPG0e39ljHvKQxzSw8+MclkwdLsg5wCChwWW5+6GTRrvuAo1QoF56dNIv9tNE
wgGvjd1pBo1LjSc3dWMgDIr+sf+AtkPmmr48R+VJ08c7b18gtkJruGno6/Jw0r35h63JTDf2cvpM
5AAHEfjCTKsDF+Ss8Duz/51pauPdx8RlJRipPdppbeSS2bvN2534DaaQWwLzdMb/eAm/h0Z+hIOG
IPaAfH/MKuCb++UqWh9kSpYFZLKBLGuxECp7EKH7E7/rg7+7aiN2hEyXPxKFmn1LQILT74zz+wNe
wFWXATjTUYnp/SPDRY4m8dhAlgPoEQb6Rdt8jvxUaRe5dv7YP7dEzdZbEN8hgHg3/MAkR4UNu7/j
mF0k3Ja0TUKVCJ68gIQENb/pEdzjLiP4zUhSK58NnHB7+WsAvyLoQg7LUOJPeqYhqFiNSonVjO/I
9W1N0buyCZ4PWNfWqgEwpZxtTpusu3pqBVVs9fRtR4s0Da5FWJ+PMP2pXvb55POjCOi059t3Jfty
jcp/KAMMxwdXIdaMjmyaZ68vqKzCy4PzzlKAOmDplT9d7kPcjaxIPbrAT8NMpdygJZmAgGuxo6Oc
ccZok//uSX7V0R+QirgO0fRcBEa9lJuXPYukWe6LPDN+kc/z9velz9I1Eigz5QFlP8/7GGvENLzg
Deh30AWfyAxXwjPyhM62Y+2CKwB0gMhXYBzJhRW/sXQVFcIUlm37t7gBddfA042zm44CtiOUfpuu
8R40yewa9xgbF4a3M9w1wcW78X/t8Xh02sQGKtSQq6DhmuMwwjshC9Jjslav1OwJd4PaAav2zWYB
HTOb17glldMyLlmtFYTSKpCN0rVDFEpQHQXkbP/quSe4lToji1Vh8fWVqkqhwBYEvyffvFFXBE6B
zQFvusIBQpfeA/WLhHGtR291GWcGNAnBQgMeKxyVJS4OA+OsfYUPNJZ5nzz7SQ3EkCBqo6wD113D
v3si69qcO0wSBLxOzMZiJB/aNYZ/MB6QV2cLnUDNk1vy1oAHkDajg8kW8QIZM6/XQglRqPgZSSyx
O6+j3rL4q6KEdM5LYopvD8du6hXhHpsKnNszVttAJ9XdLyDFTMA5TLkaEXH1MTX5CIWvbQ7SkcGR
O5Bq/SQ8PTQS80sQQByJPl18BJpFdkg31TnvwsR4jS7NwDC2zya6mfpr8Z9HbQA8fJ9ivJWATbaG
LuSjJSQMSyok7wGF2yMmnKWhD/I4xBr/B0vY+5lhmFy7faTGdX7CwCP9eNXv0ieB9Co3ne9kPrdr
bOse30OIvDTzf3k4fJ2z/Hp0VZy0gEdi1SVbTH/+jP9UKdcGNwctIxlyY51W7U6C7w9lV+KhDkMJ
yM/EA9Qu+GLeSGpsMrsYLWoH2PKV4/RJEbpjqS2MaWz4rZphYGCN3rQBSOpRhjkUBnaWFtz8W5aV
+1s8GrDKDVfbFj8629JnxmqiinLB1sZ7ZNMss3nKoH/ncb5NZdJTzuwB1Elq15TJEiIv5s5BeKCI
uscDx/ZJgn1dPjegsg507VYY12IKCyK6//UAFv/fV5obtSQtUZXPiBXRHk3n1adNc7wUdGY8Euq2
4RvcjKVBprJ1OTbKF1kjHSkTPHgNRSo7rpwzg8krVtdk+76SiqIZv4I3ygUGEGIiauo4UQJQz/JX
MH4JRhw58rtjcCGESjz7rsUxez7YvAUX+JhKoBxItykA8s3IrZsQgw9x2k7h+uHCZnzqr54kXIg9
HziXf25Jiqr1ia6yY90BBbvOaPDv3GzGnVhCU8aElHyAg/TNWA17uFn32qS9xbXKM/27py6F8Yng
01sBoyUFOQO7VRb5zCXomp2GUeg3zn0AWG1rpMaWo1T4OWdRUjo7PoLmQybYWQB1E6pMlLISkrPd
49n20adk8+0/6p9DHPz5zgXTl1FlIjmZ8vEC77lQKT/uFn9X7DdYJ3aT3RYigF/SNp9R/kYp1k70
1SpccUnsZLSc2bY9TzlPIgrP1EhqlsTNWRoy2ojWhShRCFfZxnyUuJ5Iwr27/jX7tpObNzelqk8j
H/PGBegltS0DHFKJPYhc6Ih/DgnZk5guSfk7WE7cTFvcjbYbBm096ZTQD+Y9fEVAQcPqNDoUrgyf
cAIDIQ9CCb0bFSvszx0fjGB8krIOR9OLzSBdPQqGhU4s+NKPUe4UsdW+iY+XgKmAdYnH0HLDb0f9
pvY0QdX5LF2e1EO9jKJlhTqbrKJirC8Y8Zle3y4ibrst7XaII66XTzzlC1DXXPehfIlm4V9jL1eW
jN5u3CG8/Pg5Nt9cEgks+owOARq+vZN2ZxLSdURMijfAhZiXZ7UZKuTwJ6WzMabzmI1Agk14OAaM
PYxKnVZN5uhJ7BM0+JZJ+Y7sYe1kYBk8cYmJvS+Q8VdsF4mS5jDKNK4WvYWPtSbLzUC0a5OQ1Eq0
vG+X3njew3zagMn9GkvhJ7Wsc1HJCEVv/179jVgEmnMn5pKduaBe6rZQDD4ARhXdDI9JVvpnlneG
78osCWIeTHjnGLTrjwa7pYyZfKuNCNVpOcpUXcIEiy/3sp3d2m38CnRbm+tSX1TC+NqYSeMlNa5e
gaQVCOw8wSRMhj7gWl45uegKc/R91PCkvNK+ZkuPhPu7hmfd/ob+7ZKDjg3K3WuuUg//3AQtxofn
fJNVD7CtsG4uUA0xJhfJaE375vcLwepGeFyK9d8pcLLzopsFNYSA1rjxuNLAdmc/s4FXj1vCNhJz
bdbnfZCdF0hW5Hz5RnnD8zNQxHawvglKxANavN4X4+1yU3tzXS8XR97/l5ZeG6MmblO1qTmMr7Hn
Sar2btvZRCY74goOG6JkkpQf5XxolTPTd3prIE3PPqekEKwhAooIozxvo/82WqTUUwppzg5EOvdt
lHLb3aKCGHPBzhNpmk/+jptk6YWirbG7uP1EtootBJ8XH4AFZVjq91jv7IPWaI9+uKyiO/i9og5S
YKNSgTvkasBFChFp6i6btnHbW+RX2U/UODXgFipbW1wzRvbZvWK08GmIOw2XyxCudVIBaVDq97EA
m8TWpgHHVEdzrVQsGkk5y/wYBJ9ytMfDZHEgifrE0epBCZlrhmMFhVkCjfYEHfuKQM7n347YIKjJ
7WaWcwbHbUSygTzsZpD5k9K3koasaEG9aFTuPf1lQNTJ0HCnZUCzHQipoRnUOjYKnw9Lvqi2zUtL
mCcSljQtoDLQLcz54Fiv9SqJStBxaX0YLysqqbUdbWJJa8lEIVCnVKF2zheIwju+O8o/ZKCbxb3N
Me7oidGqzJZQaZu2BEBWNdBI/JuADk1LTfQNFlkkRHJK3u7tyZgpEitr+FppPdayz4xtD+GcFXqs
6kMXbh2YIitwhEH7MlZ7949WCZGu8q0RHIulRwwdzl6donKFlvQ9oSFGj4vnmcZQNyzqhWD48uDx
auRvuOr8HMC1K7P67JmNtfcDhshb2izFrUfSa8X/whOZDW4BMcaoFKAjVIqeeKypw0W7zLJMarYn
hRsMUbXVT1w/mGiCapbz3YOp126DW+kRjAZWQxm0PyONjedMVqmzOlG/i+7zQWQZyp9qmYN/M63I
44PdluGE0KG05NYdy0y8yQtXHu3X9FboLdG2Il253zlMMY5g0No7lzTAmaoFF+SrxAyZMZVAqTVp
1+xA4iz91rYZF75h0mp1Lgez/xMOueimGdwZ4h43WmUorgosPa75r8j9Hj8uGb503BUsRyArK7Su
Fvuaod77CPit2RnRfvs3GjzFdIdmJiyJpVwfEzn7uPC/vubTPHvXVBEoQBetnCH89Oz2pzo2iSPJ
7DWmd+TiPseUDhKCokl3bEMf5z0ud4hbFaEfvPtSiEof+hq8aqlU/tydeCUutznZpd3sSYQmr8An
Lhg9tiRTDROFAA6rhEK5qPNNePNqT7KKHyaxgUch6iUv6BllGnwbDEU27+G7CdRK+LmR7fF4edZi
xO4NzZ2paDyY1mBnxc4rbU9E1OtOt3vpJiiknrshJdxMZEBjI3ZTdZ8xaqN1fum9uCd4diEdYtdb
eY2B+F1fs8QTkpyz8Q2mwtUzGkC28o6LHU2oXxd+3CHKghQC0ZqNPcFdUuOMrMqkLvQ7iltYxfFv
ZJEANgVIttJCZ8pM2KENUrgS39fKZ/lI/QNubeUmqeA1JCc6gwuTJMNsDJAvRRE9HbyxkwM1QucV
bfb1WCV9isaA5DSffHlhY+9gcH0aEBQ5R3UFG/820JEzDWt853s0HLVJKHYq2tGIWSMb3yYBPMWW
JkSJfI202ePnwoP0OxQQ4vIdmzuBfeB0UR8ebaatQkoX5iRyJrkfveL1CllDdwuE2zp1d8FOoNAl
ehwRFxFspGuH97Sx0t7MZQzJ8FL4gg5pr9Ur40b+iRJS15Hpk7qcEeq8toCIm7Z+NhbfTfycMYu0
8+R8AQn9ircy+m/rj6VZw3uMmaN4zxfQqIjMWKDLZcBzwKb6cXOMlJwDulopoYR3D1P/dFt65f0H
2JPPznohpiH0sTwW3SWcsGu6ho5s9CBom9BOkb/CIf0ZB1GLmPi9KZJe01In4U3j3rIRCvsXBxlE
+8YROb2bske5e751YfQvChk5xA9Z4qzBfJUYTeg2UQs3+TAvkIpNikK2A0xn4F1sk/YrYFzxKiZS
ZjRMYOEWNEQrzDNeJ6+906oKI4YAePnNOE5+LEfYhLeMWg5zfOFtEHcDDIE+FMAQsvceVyLq4Ryl
U1jjwyWUH/EgRpXrlLDDzKE7Gm8AGz8MYb4kbI1GbMequuDumxkXWCmf//wW6KP77WZ1iC/BVySg
C0ynLvCdRj9QEoniJiqGfy0l5aS2HpITTRcLPEe84/qAbEqeE0mfKbgrJqP8XhOpQkWLK1Abhmqc
wLtymtV1aEujmi1Zo+dMsGdi68sdSS98FvfIbu+fL1l3y1YUhZtE/xrLHd2vhrMbJhnMWnb1qi94
kfDjvE9+ckRGwSt2VL7DlyMPGt2duSuLVnQkSXMjvUxy3tkTo8b5cc9h6EBulGmL7l9wkNpzzdIt
ghECrlotkXfPWaNK7EkUTNjVuleTxesDxAR267K0J00wkGur9Ab8NWqX2ClzV8FzcAly+V+Vs3Ky
w3AdLrlXmkUYczpiXin3A1/SPqOxmY8vo/O5WoI5/SKO1MkQJOoTucLbYStzRyIh22Ybwm3NBK46
ADB4m3U8VOKDkxGEZQ7IKcxTXSi6ECpo2ovtaFurQdf5XrN7os2D/qzCBZqy3QQj4EtEw+GUGb6u
yxq/UEhW01QFf+CPiMzN0vEemCzGSaIz4N+qjZIFTOBmUF/jaz20clqyedrZtdLHO/0A1HClbHvD
qqoEGdzUvoHkGfYLbJtDDj5dHgunHNUw040U9EumWrrCek03vTHLqpLH948NSHzZauhYY3wevTqB
U4/ER3uTeQnqYhf+/vqPOIKcof9MdnVozPRgmZpTW3YbtBya712Zb76AZMUSmU3YV+7c7d/fSAFC
FsXcjIZlJgFw5+kqx21JdYLXJNKmhKHnPKaBdBUxdz2VdiiDeEQppMsZPO6kDotX6IZD+Z4/ck2w
UNxK70EJOWUNVKQN5Q5iSgPs+XONJe+83GwOEvddK2Di6lORJbA40zczEQjE8KevzonQ3SQR/l0v
j9NAHnJ7Hy7Ae8YXpPHSu2wHl53U5iTTsHFxR8qcSEnC0x1VqjT5g2yiiJXmtNRLxrXLRQqRiiKU
A1eN6SbBhbwDM8RGd1gY10hZtXevuO8SsTUsMPNuEak45EhJ1pJUgkF5kjK/NP05TE6hqfj3dVKl
2wjzhLqOU/9rMDEAurMDiXW1y5qy9VHGyCkmJb3ylPwdtbwiwZO/yyBSonGBysNLDCFtUL6Uz382
HFZVLLQe/Yc6rSr5kkkCyOUo7nixZVcjSlxLh9WoVknrWtcIkhDX1wC5ueKMlUIN08mhQbt8el5t
ty3Hzre7PpE7/pqOSMxpC7LNjcVtvBYKqFrpxWK80igT1YF0T2pu8wCvlBIigDqPBofrr+9P4MWA
H7mCOc6k/lXIIuHe2dlM21R3GibrrxpnyRjohuLgCMgNNy5u9eDo8xyfJghgBbBE3IGOZCb5wdPF
tXjvfQFRUHcF0xYxIhkGLkk8le0Vee1WZFQbQWNSvoqVhEGII1VflWjGLu2BEMORo7sr5qrWIqZg
YZGEF7RuTVtoJi/xsy+tL7ugdYrOs23qfr0GZ4mfUECfDxizd0fSYd4NzPgICjn7VLa4Uolq7o79
9kGqDDr2yZJAwNowjhU+hMMicvlc/NKPlI9Sg5QwZx4f7JGTGO5gIkMYDlxcSgP0RSZQQDZiBXgm
JSua+VllQ1SSWNae0qfwBIT2GvwBLL9TiZjmu1oAWfS/v9GHR1p8v2fUZcdYLEmHc+bMe3ibylnr
wheoe8AR37sXJvlv6XFlpxnuTNCfBRWmXusgtSR+PCHIPz/9TmbIiA8o2GdglxqXaENoMK7lj+eZ
8WWv44SbcsYQEkaKkbarfm2GiGdCqwxai1genfNBl+mGBNFC8xX5DBqosnvSgj2BiNly+jpfcNf+
FByHOOP2ODjk/U+qnHQMr+m87KSjYWx0OzQJpJVC29eGnX74+5OUyAmD2cSP1SlgHYEcvLeG35Kh
Tyl0VcqK1OVwzBRY/h1BynDJgYA+Dfk1k5vHw9HJIeVUoX8CutBox/SRgf5ONZDT0zzaDhecy/i7
kak+kDRiBCRjvkH4yQ84zsArF8cJaQKBvtyFQt21PtdRWjfMNrQgKUvn3wXbI2SvhJ3RYwn7bfRC
prIlLns0CJLBPUACNEqXFQ2aO20fUKGcstpKh4VQjIcK6zGxfvXxZYAyG5NRlwcxpGNR2YaMrmQ3
Lw0pSI517R1ewK2OXZ4HgShQu2AWN6pGlOJUBhmxTyMd0KQ9rZdxGvjybV/afEQVmlVr7xPtzCVW
CTxMpDFEVWUeOPJaTUs5tctmS6Ecl773Nhg+ZZZ3STq3a7zx+lQS0fOoCE8pHWt9g7/xjI6d/hab
Hwnd45Dn54OXWw2zNraIz51+FD1QSbl7zaLrzSJk9qWUsRxsUKXAcdkHY9Vq4fqL4r80WLszgz8x
Rktb49sCbgvkt3tANlX9yjWhyeyZ8xoHGo2LgCkUUJnZCSun6eapEy/A64FFK88Q88dkvSOPRkLt
9lD01bnHuc62jfq8HQ7TSvquStFlPhtjHaCGLnARl12P6ikASUIz/hsdBJjYi/m/p/0JP0Varx11
G8Bk4+We3FrnCGxib9Uvssereg4CZpiJBFUdZg3Xy0ingLmzVP9RVE7NhfCWpe7NWt1gUk7Exaee
pWcdKdw+F9xICSSCA5Ck9lIyRKCJwki2O2xZGiU3avBsPqoPCaGitsnxFcZ3us9Ld95zp/TYjjap
mPNFxyWIlnF+77gzoME3+UjQ7GO//bEECQeSNVoSiIFgVVpgQB2ZBYoBZuJIIckFEYnbe+dOOz7T
ZQe3BF/XmfiRIQU+U4WGFqOqLM8jWRiJ+y+CYJdVZoKjx2LbGk0CoJsNrdQ/v/qaX12EiLjhT6xs
GdJctEzaiEVyLh+KHvZ6M4EhwNp3VX93okU/hcNK/mHkKx1z+2TxM5x8qhns/I31kHzb98pg8xK6
ov1sGf6XNegpbD4R+arG4MuRE/zYtcaZiuERr/QeWauImcWKpwZsrP6k80RB1su4bvS8jHezkvHz
j9x+RFJhsfFu9Jluo5vmQjjBege+E/XNil4rgvPOTiabUbaTSsaoYWpzMuTHLs1zBAQKCy0Qd7eN
MBzXeQLMJK0zwFceOH5JG380+NHXeFrreiJldeROCIdd4KGXAYSa0ryDLFilsYvFNFW+FQycwwJB
0SssikW7RVK3yWRTD5eA1nqltxGHZYis9c8rplwdCyXfThdzYMkIgXjoy7Ct4MdFKeHM3Yf2w7dT
yeB9sBZhfVwi8W31z+neu5Fh0Hvs5F+s39daR2rEsugj9ZhLDH7ovJFsU/RvEZxmi4it7EJ55Xq8
yb4F92rtAO8Ve2l6ZewkLU0D2U9jgXxX+TaGz5ZNZESD7hzGOQfE0yoIgNmytXjlpYMbV46qedIH
nYWeTIL9DSFlE31j7BRmgcUv+IejMW4G0PzGQWLwD+1S73u/IdEejZw2p8OTcQlI9SFMSa9FjjrP
57wb85qGuUuyqaYt1Q/zbN+DBKZ+iDVC+dU4Z/qPN9pIZKHd1QX35KJlWFsUKHKDc1trJysKJu2l
WZH3pUoDLRe0WSw0RtC5JRXX5e6+y4/XC/bR6iRaNlHRAtimX7i/mvDUZXDWlNGgAYJpp81sTW9q
y8yE+6mCzfpbS4fEGJ57XW3n050Jl2JoRti5hbvnSNlwc1eJ01aomG+VJWfHrODPfsG+PHk3fVul
DBVJKw0wHZUeo49fHb4T74ErVEXOAYXm/KQXT0r+U+04R+dj+/qELXWWdM78tOHHq9NF1x5Ym8zB
qDvThY1EoiLs3Szj2LbdZdxebqGnPy4eda73VI0t6RHoZSRgrqtiTWYM5QvOG6zNyeo5DXRd9dQw
vQd7ui2u9KXAm4aE5cVDQBHHdFwalsGUnAEWuJp5F/bxFVVymQpDW4hsaAAyKlL8615tCZXYpKp7
nTDl7Ak1r1OM3wSYfXkHPdxlUE6aKyxoLQ/k8JGv9sNqDjJAWpoKvlnSHP6ozrnwYMn4FwKLYq/F
cCOFS7YXOC/ypRibjc+H/V37bir/xXyXBlSEWAUq4sruDy1zQT9c9bLsAs5ArYJgraKvVmgl55NF
xKndABKHu9vMNQun6q4X82x95qcpBBJVBf++TsGXE/fq3i9PxyGP7mWMm+o4FHfD9H/W1l1RwR6Y
6Xe8+TShc4xDL74S2aTtovtGsSaPbkjBDgESobqR9aUZVsw7gdMpwktWfAsmxTvbA1CdXEpjvqsz
xjhixz4LJDCD8JOvwXgat5HWneGTlTNDYLKquF94xU4j/lyKf1wuxSF+PKR8eKshEjucOwuekx6A
PniEkduxCeHVQsUuldEKzmBhFkddG3TSzFllzCZEJtMKGPPXGL8LoH8Lj1N0uUPNu9n9gUY6Yap3
e8+GOhsmrHTae03gGXmjFJ/ateNrKhE0WemEPq+GHVaxw2ExDhp6OfEWHJYftx37DjsWiddv4GPv
XYhKzlNYAz1M9GLFuHHMUBLDba/Z1u9tZ9i2HyI8CT4KoRbn4m/aMTLoHBefT88oGA+VB1ItWT6n
IZnUwAEDPh2ZMRgyCb+KzKIPAVcD1458GveJcO08yEZsyA6HkWIc04XgS+zOfQ/1mQOenFY3ESRj
FYh0UY0ot4TNsZQLCNR1Ks5u3xsg4IMOvCFjOFMFzcBIna+7U4n19dh0HdHPRyTfrvUAzF484Fyp
rMgIy+k6GUu4Byb6CcyFWpr1nGZE2Duem30u6EWTFYwbK0e06tIP2DnmwtoRZG371Ii9RtXvRaNh
lIvxdjhRCenPYjcOLkaDzYEcBeCSSuBX/V5btnplQsilN+Jap+x/V2YFEhDytRlw6a5mSS9I+9Z9
GiwU/+NCil0dgW4fiGiO2BDo2q+UWtBZn97jSJxwIY1pSXObJ6Ve7eAHc7A3YCxhk8EjpCB4nEnL
RPrrFJkDzNipu6Bj2vewqt63Cq2oq53KkE/CBToOVym6uPq3k0D+cOzsCuQ+XliqOBkMCviqCjU4
uRoKoESWnmbB/GAB322+7qMKJnbV1OqfeiOvJnM99RA+wQs0ClNTIMTtlS0NwcQE/vXuSPBjrwWR
nkfxJ8MEaywP2PQG6EZ5QkG3rOOM3a28DzJSa1xUJaP5OQk1X7gc0jB76uW7T3FtHp3m9DkB39Ul
06XBnjal1OvtqpF3Y4jvDrJSeb/BZZ1qD/NZm5qZBb1ZhkggZ4ef/La0ya1hNJVG/Oyuof34SzLt
cy1Nlmqwzzt1Mt0iX4bRHSRE76YQDzRvZaJEWEavYoy4fuMpXwzgxnw68Dk2OysEhUipdeOu1wpi
/dj1k43CO6GdgCWjWVUh/y6cG+6b7Cp8VJUASlhez8tK360cKm5rNRzcgz2qbtfahaiI0QmJzDuR
iZrc0LZ4/yvJwP2IOwOk1orKwuR7nn9XfXEy2nNZWgq1VrPoeaFTR33lxByQ77ooji5VUrGSyGIU
02f0mMX1K1AJnq9JOrphC/9aiyIcmo6Vc10gJB9QtDrtBkCpAKxf6YB/Ej4mf1MyakQc4k2Nxw10
K0AvY8h7wqrhwxOknNvZ9gtREH1MOFh9sCI1oC9xsmvzWPcGhSMOZH//qRs67ybtoAPlEHnP0Yl7
hOSX+NgVtSzNJQTH80WshMwTlcSSqHDmfwqqjzxryQ8BQ8+ecAjmP6fdnKWaCsKpOy2WiJam64o4
xKq4C8n6owoeYZMtzZngUMu3ucBe/B1iC0xlQo7DdXmH6URZlirSN+w902jlbOJFQs8GnVUID/Ua
+zQbEUxE7lpOf0dUz7opeRenKuODFRCL1ztfkrDKHGL0hQixQBdxwyphEV/ojXUbFobqdkvDyOdS
5GsdrDYA51tbPt3lVSdqSxeFt2p5zMH12pyLp/Vd6GkZ77lvl+nZBM9iI/nZhrf4RJVUV7YXhsiN
AZMFRxOxNEkCouA9RH4dI1JkgTzLHD3WZlBwXsdYZmiJGi15SsdxJEjmKiKh21GInfsMcSJjqRfM
N9jyY1r0wgNA91eDt9xWP7EtpGW80Nk0tY/TSQ2UURiV+7VKPGAlePtDv+QzUjVYUSGDZL9cv/2l
jSXgi/pgkBCZ6cmGwd7LO6dzJtyxwlB4AjVHcElFpQaagQQJnuR69iexiEgo9YKNeynv2RJAabqe
GfVMVJx51rtQZLgSvrIJUf5B+Cs0qdy2hOWR13WyBLzNgxbbmae1UTdvbeG41MdwgBQvQQej3UWj
QbkdD4NZuMAKSET+WTF+LgJXx24hDY1EuFIJeUEQI2NtasRBh7nnjD4KKNyMCVJsD14zztTK+DA6
3yx2QZXYGkAupdApYg4LZVDDziodbWFDQyO4amfD2D/6M4HZ8+hQS/gxDFCrn4ui1BfOXmGT1aYT
vwEn4XH/kf9+RsQPj0lCU5r6sbXxxgBqZUdnfZ51epZKcU3lV+HKKjT2Nr5pSm1H3QKdATxJQ7M8
t/vuJuuuxRNuYAkaOyzXfi0IyG3ZeB7cEC9MS1RyfI2NgLBPI8APwCsZhzBm0PlJSOwLtljT8a/u
cDsWxstmAoTZvHL/hzLR/eIGkWlqo8u12eaGkga5PvHelfVS82xtMtw3dMQPGFgyuXk+8CNwsruw
ztrWBvKKOph5a7r7mcCVWvJbvJbaOhyIH1dqzGAeonrnuer8sgokEpZpsxYN/oLr/So1sa6fWncn
tKxBGzapfeS1bLBpubdjfBgLg5M6przpMgAwv3EMpQz6AZbfdVwA4zLH4t7As25AnZZaX7Fd6AmJ
zr1k1t/3OP+akCC66Fp2mlDka7w6gQlmCku8Ww3TqC25naOxFfJyGJi03Ihx0YG8BDo55d4GZb4V
N7QkZhkFl804GsLR0Wsez/5cKkDQN4asns3PAgBufg74u2xadWFIwXtrOepU+saO/Jx+WhWm/ABz
grfAxsOr04qhXKBO5vjDBXNkaMDL1OAbEgPn4eJNqDafyIaW+2h37ESfFrMQOYgMB66rS1bzcrSO
sdhtkMgjDbhtuL0DYdSPlgZNjZRnCumMGmoSY2k9bjLldBV5iZ7vMYHldQGWv9UXC/mIZ6wHZstd
o6zaEqNO+ZbD19ealp4/KzxF8WVjJ0JoMkBLUxlXCR3yHh17aRiDm+IVUijS5aAy9ZcWjzK0oKed
HlboZKCiwRvQ39VgqHVXYyLcaWsN7B6g6I4zFlbjlvXDbLSDwfbz7hYiyy1anFbwEyHzUuQ3uM5L
TtESiH3UGia8c9hbNSqcESIsdEvxLk83sfTegR9vQAJ5ceOQRKJ9sH8vzQ6kwf10BWLrXf0UCWuO
lrncwu09JNguQ2M6P5CiymqKNR+NyNTmAhIlt8NJ58s4aQRYNgzOjNlOT3pnUvjT+wM1rbiqtdtq
h/Db6/m5y3p3af41fdNUl3SDT9MrgLg3mHyF5KjFU6rGQuGL9WkOyzqMsL4423LKwYz8K6UlDEsq
kNhEIk/n9a8zO/UdIYpTCw6ocCQPuxaAL0TNtcipXfftSpaOnSxqt0PombEIARJyfOWOiJCcyLQV
FV/HxCiFDER4jmApLayX+gmQbSNx00xgImd2h4JDRXz7qTVTStHHQNN+1j0kU00rQnP1mGNSq/3s
6QTC64xC8Z/cUeQ4I8k2o0EY7D+j2IqCPBnrQ79pTcnjjk3aFUetk+swyrk5zE6c+BAB2S0fqrQf
Lina2Jpsw5dr8jMmrQEAb5/A1KwlCmfhuyjK1nKJKg/KrpTToZnYfpYJ9ht7l454RuvahzocDVI2
yo5iNhYR/ruT8Cne9yr9E2O56yRMyEU/IKjdHLcz7chV9K3W1M5qRSsy9eFZg6CWCO4vrJEIxwXF
NXAfOTzhdx1F/GevmAUlCkXMbLt6vY17T6n0O6MKRFMt9kkC5h0bdLXZ2S5JV2NLqtrlQkUWT7/d
eFqAXN+zSMd/fUdhDmPV5AJY5mH3cHSq1aTDO/9sTvLppPbbG4plTK7etSxdNxtAhATSjLKaBX0T
pKZb5G6oyYIgCbvI2iizX1wdpOyOis1ww0TVwHXELe6L2EZOV90n0uD53uHXwvycqtURipmlH7je
6htCZvYOsOaVzHzTetqCtizRktHsyhfEjBVyptWYjZRZzeUuFRGfhJeT6UFKYkEr6mqa8e7SmYzy
yTyWfo/0dBWiOqdQQWM2wc/0eAolUkYywB01DOIyM1XA1aTUmsubiPuUY1kagsjrVuGHt9cStjVo
8eSPbFKL3dKdAmT387UKx/Z6pNNW5YTahNHGKQWeTW0gxXam0Jiv2enorm75Ff9Gt7Dtq7TobP9h
kY1XUhabcs3VUWPBiU/bpFYcfDJ+J9KeNdBgim2qgjukC1QaXf+NT+Hxvj7iKqk5zRUqunz2fXrw
5wAL3eEWdHsGEWKcTgPxU1CGmOXOLhRNUzTVNyyGRMhL4LEAUsxjhcPuTsZRM/PzN7bp4xo70V2C
YZPdkg+1amf7nXoIWgv6LNUdp+LyTjL8QT2szvBMd1eYTQh6uj9SxUVkSsgCm3ZOCg+78KKjP4uR
c6ZcY95KissbVjciJnhId8g87aiXw9NQVKSeGZ9iKMqf9XvBVzKrljmux/ym5k/Z8ynre/m7M8hb
kNDaw0LPes0oISuP9W2YCSz1FZALKTlD67XnVEuP3ud8plVUzspH2GUaSSSZSuJpruIIO7UKLG08
EjKxzBVjophWBJDHFUVlSkFsRfsOCiV3mcRFKO6KHt2Ayk4jEXsTVxTtGAn6oOZ0uu65eqZTEvuH
H9KqXUGgVL9t2qzG8rLkWrV+QpklrejhqeTbdLtCV95LF9bYURGvS+bdMyn/rYHrzV8Xc9T9Xd2T
al8SvsxuF9Mmb+r2Ju9RvSxjTyuSxWVdbVSQ9zR+PKkhAtFr6Joj7nP4Qds4h1etjGSEG10llHtG
I9JyADqTBV0skmIsWcG4hIInwzawiOf2a8FWQJ6TvUGx/WYCF1zsJLPTrmA8h4cc1aci9Y1RgsKC
zV0rHGHh+g3XkbQBwRE2jkLMsEWOwgSs7WvajjALr9N6qHymnPd/VcMJngdOCqJQLn6IuBaDhSHn
Wfo4jrh93gW2Jp45VU6WmgMBEu14wNwwZVRH42EZemCOkIJN0fEUMCw50Z79EPsxXr1060B+9xST
3rdjurNEJRimnlhsDehx8cDn8BIIlqel1vpxOhDU7pPbY/KsygMtudewhZ5fv7HG5uxdQVdyBwIn
12+xRpdQJYQ8T+f/45noyrd/EBxMY7URLHgCEx+SzRW29dkxffkeELigJlmp3pmXlxwgFeRnYr/m
gUSP6PAoURicKX4OxTLKU3XfCdG69FcMbdwxNxhy9uasDPcj77bxr1Z9/cD+MTIAs7qaXhl2PJ7n
7B5/EJbOWgD6HH2Y49br3U+f7ha1nerMUBn+8bSjeca2BlopSKyqbhZecPlLkHM0X9i182vNRiRe
HoYMDqY9SH29kwsAqz3QAFO8Qa0ku/78oHUXJ7TAEnZ5UHLIbAecbFdvVvrzPOh7X8g8hfnYe4x1
QGgsAiiXiKfMpSn8dUAs94Vt1Zeb+Avntqqg3JcJFLWIpZKeSlvO7U+vmNL9O8EUWvtFd2wEYKrP
nJ6jGx2OvVg7IeVl6RdbKvc9FwmYIyCSxUxpLmWZmK5lWCJUgq3K1iC9clRbICjrexXJcvrW2K/m
Mep8gLH9dzq8qriZ8+N7da3TZRK/4rgMIiFl+aDis3NI8lNxIIhZvjiH/Arliej/XEF29m3OvgHC
TEf7Xsouksjbo/AC86VNFre31LFM3npgZ9L2G/QEnAcB/LstYYOWNhZkVCDH80BWEFLL+mgqx9ka
SS45ERGwWnPa3Djl16TCvrV0zKSRvBBlnzezv/iQcDKGF9s1tYomMYzSQmR7c0RxyWiPNCp+hgyx
RMP86DrJ9BbByG8z4gnDOBfM2usAWj8awW1biANtYfVlTJTTI5cnpGr5d6CeAj6L9tRQjBX+JhdS
K0rHyTHj7METFAU6VW2g0RjcWLmkatRo6pDwVXUaOEctCbRLpwER1ZIUU46TkCpfhoxBPpZyDN3B
0KBH0wcMCE0mIEbNgCdXv9a63JQia/GxukVLYdmXq5UOTlPmoBeiCFry5lyPuU79ownGpLreZMBk
mpjIxmBx08MEetP/eqbhtM3Z3qJd4agPojROpy7Ik4TrdGKMtGnPT/HLNbdJutnAAx46qn79qQRo
71fBu4/OTV+bSWwpU/dxOR4U4BxpRezDKCqPkTDcL4shiy51mufMbAWOFTyK4iFvLwD0wXkN9L48
xlGb4LeCjgV0OIn5McFjFig+QO/rBBsKYdHIpUFapBPBApKXquTwGt0Qq5DVBiPmAdfejnsO8pKz
61q/t+kc95gl/3ig1nhUpGIzxj8S2yUZkjcUvcBfIaCSukSUHzPNlQM3yc3CBkv1xrIOCc0J3OTD
5J8bhhFvSH5YByaL3xxwn+klaAxjcGPDoclt77lJq5mjEMaR26kLdgOcKF52EmlUubiZcvuLpB/H
uE5WMCNRIBug0AaOxGU94PgH6//kdMhGzY+yDTmGKib7TYLvjVm7uePbDj3sjQuVkfqJg03yOa7d
LO6hokVTJ4n8uxhrM1bVgx6NAe5rnvle7Zkq7C1jmeNLv/5fTJozXoBD4GBAo99RI9REChNLkSQh
tt18szVFdohQcWVYY8/gTV8KfcIfx3nOW4yeBK5TdX5K79hFpFFGZWmYN9t6cfBoIj61oOGc0wXn
2WcZWCFqxhukCVLgYwgNQbBoEiqMarAGAB6NTGXg+Ebf1w35AH0IcCUGXGqHQXoOUAEzHpZqAVsn
5IXbqkpvIGWAeogmwR+xz5BG/IWnHodctk6tJcQooM3H605L0S7m+s4hAvZyTEen/CgXxzk7Y3C5
QU4iUuSdmD6jtqOM3NCvzRtiXpHr6D0IxoO6csVsdTmeipT37Mygpwb9/YMuA7Z9SyiCrjZ64Zeb
iRhr/PWtEhOSuEQmGvUHlGxJxsoWZHmjwciOAmcjSrok2uKoZGxJw+tn+fuq/4U6UI0yR2cWuRFf
77uX9r9Xj18kUqE5NJGGqpuYu/4mE0+O+PQY02yX06ktKGXq0vzsGagInUzYFKdBYvDsdnXiJ4f7
CF4AYrAiMk31p2X8RnOqx/VPOJhFLJjR6w01R/RpfZJDV3xiIF9oJUGNnjor1mTGDtsREZWh9Z7e
ezpiFkwp26/5Bs+2oD7tyrqGWV6DUObcTII8MgGuEZyhc7QEUmLZ/END0IJHOQTBX1MSH6TaDlId
mwu1lVGly/TPeSzwZowLlT4L+fOMCM+k38kdTaWX3tgZMd8WpxTc8soCDBf0DJF6yBCsI7e6/AOK
LlPDAzcI96PB2cXsQRn0Xl2CFsTQc37emhvh7yWqPDIuDg7GVRebVkuXg3FxTu4aOKUODi9BdVUD
n8WC51od/v0M4rpkSkt4cgBoVy7pvMNhRslUVkc1bQH+jqDMU2WoDY9fW7d9jrNmu/mKq1255y37
+xU6u6+28dKBQkuLG+pbtb1m2WVr6w8VSeVBiDfNFhlIP1MI55L/xp11fHtGDbQdwdnntr9Pou8m
mzIlSn3yk2vaoVWGO80ng+QarTwxIryXH66X2dvqBHoUPLOCsuQqY6bYdarFtsSI4OwQvBIiCoDz
2Z61iHCPQa/AYr4LZNmF05NGZh6JjRg8wDVPqKhqR+AxpQpedue5bZ3R4p2b8cOc5z4OqHxsS2KL
cfvZF1WIEab2xFCXm+KOZ6pJq0+i4Dewe/BWNWU2uUnSeLYy33GUdM71C8JB7b6uL8RvjJjqKGWn
BVboYIfg/clRY8cy6tpY8B7+TLkguJnqOJyKzkm+rS6GCc0DmUrAzIjAnO9Utahsn3YLN+MuQ9Mx
v8L+NAphvReLETtD4nFkAjSt0Z+j3aqEmeBEdQrBKZ4N59iMfQazf0jMODhV6ZE+jWOINAaBNdIk
uXPwLyxARzZQrXMtDTpZrlKn+n8oOiFBZTfeDC67mLa5yNpUkjY5KfsZgjT4vgEIsjzbPe1lGwkz
FNscIUcRKTWyuO9wLcnnGW/WmuJjGrwlk9w7vA51TnH9HdRF+dja8xfGZB+v3cPZ1YIVodb9tabJ
pfwKK3hA3iVU7ltiuPsB8muJdhU5P9nO+p48kRtNG7zvsuYZOLnhE4yQvzZTsoKZiud/zEG4jLGz
uwSPiHp1f8NqPJRXqAe5oHgBVjYhZ7VvNWyZtZFR4r16U23/zTaXsTYMqTqH3rUkdWBiLCZFnUzf
MoLm5MsTn13mEe6H1EabVzXCy3Ef4sQQfoFXX703hzrFSWi6zpdE/gequ2WnrieWGiqXZss/rji4
eQyJYrap9PuiKq2nNMsi9+5XcvjME9w9dMgmIuhdTHev/PXZRZDRyxRT9U00y3UHczTPcX2FALh7
Uyw82QGFtrOJhk2BmmWGZXOng3VO+htlA2thfhEff8hMQxKoc4OMUz/Bkk/Z0EZ7DkfPZCC0QqrO
nAb6AH5JH28N1bOokr0aXDbXOWz7Fwg6erw5kxdO/MG7SfZg0uKQ8f68dQYDPdeZKK8KonvBlfU7
gBrSsHWSct2mHjzRLR27693Ot9LZLF78iFqUGR4XxdKWYYxoEvS6C0X0ATIphsFQwaVfFGtOnITQ
PZMD+eJ8EMgMpQHjsY7YQD53bhUoqKObTG0F7Y7A/1B+KwYSREVVKdjtebJyF+/8mS8HFHoDohfk
t8zkZWIichwpYGGpbi5QrXyShZGWmDHv5Z9RcmVYP9+rHDlN4jpsajQ6c0G0osetAyDf9ZTX5QBf
WWLNA/v7OwAy4+MAEz2L3WolbI7YZQxkWT9AC6C7FCkFerV/qphnQuwsN+XduGT9n1S3jiC1YbYY
GeCCHlNH5ESzw7HL81tjy6X5aysuwAJjkkH8wbq8JIVevXpJlKdfyCKHdAnzY3cdRPJeRPWq06l5
EvO8Zv5o4tyjOOBbSnZwJvTp/q4Rr5WxAmkjoVts8x49jgzvd3OdIBfo6eHo0DRmC/mgK8i8Tab9
U1SKS1lxSWoCrui++qjto488WSKJtELSys6OnUllbQ5H81fKzP4hlZGDWkWN+7IzIYgBoeHLFRQa
liTxSRgJg4ggp3WUvhCpJE4Uz76qVGzgazr8ZoXz9RgTpqSuGAHrSFL8uofCHOrWqyLD7k3tcStF
HbzKdQNm3kaH+NSnCLtHeph8klgcEcPE6ZFimv5kV9A5pUWJTHJt9dVtL7QM1hXehob/vaj/RWql
YAKGLSOMQjs3acl0geFI3SpqAU8tLX3xyfoS+Ouaa7VBMblQiKNkQBf/+nYvm1LLYE6stTBuTIcU
cxIO4m3AUJ9arXY5AQa5xY/tC86cLoDvdpE0zntOg9/DgghvKGd7u96t4XMUvDP1oKf2pBeFfbg2
EdsgDNw3AaUbVAPgc2NNBQX+S275JmQQYPZHtdG5o5VhCR43vBIxdTMBuejaYSfveIIYZli/olgu
GjpUepVJmK5GdQDnrr3Tij0ASf0AXVFe7Fr7iVDCmyAnpUeiOjpLVtLU5Orufba4kdCOwXxN0S0X
Pi/uyLOm64O+S/1lQ6IisXiJ1YorobEvombJHYsF7VLcoy296FTATJg8WRnvXP6Do5hYL9p/FTaw
3M88L1czFqj6MypBR8lPh7OQOJwgNoEPgizCGznrIozMJSASDm9ysWb/SH32OCcpTvPetWni9aen
DDEhHZ2w94OBSoZKy4pVvMWU1oXB6RL3Y+X5Mzt+9aiiXRPZbn9ZugDDiqxcTzrxk/c6axCNmJRN
4sRjTuM6FfHxs8Y/SHFsBgRIqIOVtMxofi/g3z+9/FLNZ5yNXote03bCQZmXyjjs2zJWMjZQsnIX
UjHCNSXdSIDDnVaq2rbBuah91FczGuNkYVa0/SZhUmPwC/KEALvAYuyvrB63BTNU2kfn3BTt5r2f
Hl9LhRUPBRk5zR+8T1xRSS34jBjSK6Z42WQrgmNUTkpGYb3EgmXmhV4xeKBah4xAlr82kCAI8LPg
/R2nOLD9dkD5CoyGNMVkDZQMNEjbLzhHmJ+n0VALCtMUgY8JAX+F+0pCeZO6zTvHVCLMxIcOBPFI
H0mMm1ul8Wa8ke/a/+hb2GZVTCpQLGONHZh+YDOL/P2ajpsadVDnJl5kxVz4kLpyUIvJC6kNZvoP
dqgx1t/+3GhGmiJvaMfS9hE6MHQkWOj9z7xPlyKjWbCnesM1m+E8m2ZzlO0zqtZHJPOHcX69/J01
+5YuE0094XIokBe6LpJ3y+LB7veunL4NzW/1A/EZs0MXbQl4Jq37nxK2fqQEdwUsH83FZjpi9IhR
t9U+ZyyqSMdG+CCqr5ge7vl4FPAAd+NNmkf6eofwrwUT4A1X+7zOsQJ/vMQh4AYCdo3jRB7NuXeF
hY/pndxyepQ6qwauqpZ9FQ9zMkvRo7lJYcm6FoxvaYpaSqpKlO3yKqBCqkIX+Wb467UE3zPHaV7c
FYQLmlmPHg9EUU+IVM9ddHD/5Mp450DF0ljztG05SnVEEXumQOxn7NyZThHXapnYYalLwDC1l88B
dxu8dVB4p6G0TVRPjM6gaeKPDkosu33fhAzCmFmKRmA+YujcRGej4eUmxywG7EafV8gVwrj1xx6K
f476Q3JIneAKbgGnvPvzjOWqqkdF0CVkilf8pk8z2Pfqob74S9kBZkwROT0oQGU9QmynjJ7TU6mj
LuLT9ACkvoJEmWf4jCNudApwCxQEF1VhQwWcLMNk6BlLAzmO0/A/E6gNQbzA9St4IyT7YEUcGxYp
VBeKCzhH75RbwKzKuVxFsIQPCmK+UWaHP0A9AiRNvMwQ/5DMwBMQ/R46fekmOz82EEn+QPr6g1/R
kCsA0oeELYwLNpA6yxhaGwxLObDOk4agy3yx/Q6XJJzsZIvgrGbvQkyYlhg7ah8BFi4EFNduFLxN
EmwjFGQoeP0C+bucJcT27rOYhprYMk5vwYxgd3F8XEU5otiVtNMSm5GckI2RNY/cLApaTnHRC+Lu
b0IBV6YPRiKTuPv5vncVTdOWOOy3wphxHaE7niMNtIEG9FsqCQ/SV2CJP4wWlpMtVwrGXCpAU6JN
EDpw8/WBJ/zEGeO/9AP/5KJ0N5mJVhe7uJbk+BqKUFgwlG74BaaRuzxXezKVD4BhzdgWHBVpU8Zw
g2vBnVjmY+n5NzLJUnqTsELDA4Vm6aCOajjUPuXmuEsAXPRpOTZPPMf+088tOLMEVg8dp4BnatCh
FnZzOzENxL4kzPhkCyNFLkZrq7SBG8Uip86Zt9Kvp56LBynEGKu3mzWa7UKIwtodT7VPZp7dBsJG
kb76AAhxJoKXxxMMw/rbNr90lsgI+PJmlZNaAT+6iWQvaS4LbVNSf+P+9rtmYfbAyEmUW3RoVRo8
aAM0x0clp2+JksQWUOCepT12Tt2FMqIuJVXX+GT1l/Bs1Yt1CpnB9qpf845s0V5KgWgZCWLo4Eua
ntLNHI6xpmzXTLZxt3wCPhqg9xFR7s0n1F4WdFXr76TT6h4QTlW8PszjXw1RCiZ1sBvB65yPQEUy
4v7jJEPwuAAwPwSc7jE89s7tQSQobUo3NKqieK73ojSyzpwA4N4Gi/PFwqffOGMtOBTcf3Wcm0VC
MFKVkbRc7HTWdOE+e+q3jGns04qVWhzmeucTRsD50X+a59QoyXyhW2T52m3JwlT5Ao+v7JL92Vyu
agr6XnmwqLjPcQ5Jub25DMJgtDjo21v7RbESS8xQdSkdd2zfpvmhBMj1kpzf5QhDfbTEaBG2KJyy
ngnBM2kRWM+HZXRfoqu0F9lhqO9+vK7ox9bR6Ds14WKzdGAm7X6oPGazFAIZzCpqxHcW0aMiSgWn
ND9C5ovfhQps5I+56a1RsT25ffcBb7BfzqRb6SNiETW8/SNyRwD0spk+zGelqP2h2GbFMGA9bnH3
DdCSNBKiAdY8Ps9Csv+bEIEYKwR7NykkbwevQgg373CBDB0o5TlpVw4k7HBw2RFdtKep8eIokP2F
gQoh2aJFIGrJIxFkc7UtVKpczSf1k2eIzF/v/epF6TGbT1WKI5qLrZnA1MeTYwNXUyph8E4RIUKW
zNvHsjOWvjUzKL/uJs/8MmrZ407qxxvxhvXe/OjrfGx4hl+UGE04xSO6QwLS4VbS4dgboCEGDSGD
O1RnYwLPbaGX8+SbC18a+2b/9LJPlrdOUjJa4wmnB/xW7WZrxaPFaP6cLUZC6VB5vd/2SMPbxYWk
HsA3r/ID7wBiaK9kugog2SgWBFrwj5wbxxZtMttUC3cRaKf+s1LG5IXbnQ4SKH+X6v58NgGYmdZ0
Up5ZXJCr2jXkkjHGFjXrWyuFT+tAR59mjoZL54R18hQHc62JuSJ2fPYfAC6ePWnZ2/3bdS8pC+rf
PzvUmiD4NHQnW87pa666U9O2abOyZa9W4uVbf89BbWD/CKxHqbHMOEdaOm42y/uyKb0vs/E/DG9v
VJtZbV/RvX0wW7he5RP/kr7PtZOHxEWkvsTKjRjthXFuPxBjFuVZ9Xs4M3QyqqYzd3FYSIMHV96G
+elWsPiObKdVRxwLHM8bStr+uKRA3fIy+d0jsunSv69U+UgnwH38iSE4+fEZkSKZTYYUSnAaJWdQ
G77HF5hELaKmgb05Cqd/zEQQ1h+9dQrfclTUyj0wHq+aoCbW6PqkFCfahwWOIFY8rYCs09Iys7Vt
qTZFR/4rMYlvDB3p8Y2sx7ySilqqdTDsFRJjrzaN06VbFw/3NJGMb1XYyqa/zuILxlIzTwp/KUbM
11bUDw4BkxX9wwhbVW58w9xAUJtP7snDDnlKQ3j+btqIQzReGP6E69tn+CY2w1QEObt36jDeEt97
cl8TuUx7UxMjIHLEd5f607k6WHfXjTxObtn1cjTwMSzrWSHSRU88GziaSv/6fh4vMqlyEIJPlsZ3
GVnVQg17CKjgFe3SSBOqWw0EaAiiRhkbyngNad4ji71DERuDWTQHxlYzGZIKskSZtENw2fbNVzL0
LvGoqgauN36BmFgFE3sFFEysmrCIUNO64fVd2NS0b3HF8FB4KWz7P2D0Xh7daEpJ4Wt1HSdM0eH2
tggy+IMmKiwoyi8iqv6Vc4bit/ugfQpN1etqNs92IoT+jrsTWVqPxdFI6zoHAE8tNJslLC33kO+C
2rgF6zOM5selQF1j/ON0zl+8xV8AMe80EYOgZOkzZaEDcb/fm2hgxzgdNAoJn90qqpHwiLpnZ5Wi
0lB32JJpGiwm99HTkba6KlUNhmHe8AQC2BwrFf1A75WssUcGqz9RLLSo+OvKJdF6C34wWEyKftHm
D/XZEYrZkH3muekP977eVw1mpT3uOzONC4oMPNu2Kk6sE5u6Q/IoGRy9JUvcBZohifhpLQMkB8s+
Nsd4HKfSHyESBBafnaW9hRUouxA0QfPguaz6EcyGcS9hpXqNrH8Daqvw799BWkPD6d4R6oIwx/8J
cT4D80fK5bqGyCtqt5oZRaMY+WkOk80eLkXyDO9UkH3e7WkDamcceXL/WtvfVw/XjOI4+ba+fMl7
8I4od5m3YKgjjNuJg2vfJLayfSHbSP0acwnS6AY3FSvXx1sPrTAYdppoJE3qNlECrrGuKmZqxQoZ
EcvUcqm4d76V1U//ZH+8oHea5qheupvPxeHnM3978ZM+Jso6r9ykmw9hXwSj8ncyjv1JaPH5xqoI
Eaugc0CvpbPQAYXqEyA3PhlJ0OC9xZkfTzUUiPMLGT1sGdoG0r+5Abg+tTAGb+9yTIO9e4SzqPct
wcX/lQLjxqd766TLfoZ1aUapUNvuHwRj7aEkyHn319FpSXm4di4RYV+GlmeZ92veAN+FWideEmv0
kPxwv8Atp39meeF5+lcZ6jRDU8Fh26cokhOulOoG6NzIY0dmUY2UM2TUhN0iUhjszbUw36u3XWZy
/TvGRjCLYH10MXaQGanCmR4pTEHPtu82FXACnpp58NGARdOBTWazUbCBXJR5KPU1pfiwlTQv6VIc
8SmHxguGLE4oWvqWPEsU6HtedItXdmRugWOOYO1nI60zK5GIjyhT4CkWLsRa7YHZDjZFaQWL6qUs
lblscVfxs1yY3F6wb34oYIq27cXD4RF8hw2PRHMACfLCJ+M+tbR6KA8oVW7FVqmP0e39MTRR6Ww+
toQMpN2Hi9I8BiVZ4UY0jQk/bD0jGU0QKSa75dZFUv/6f2N4GdPYA7GyN/AZa4zLeMDFH03toJuD
h5wPm8kYDIqujrFiGgojldlegevvNznVmEDDrG19lGkiR9q3mJpBdVx/0AWbsGjulFeU3HG/4Rgx
rc1o/olRJm8TERNdR8EYOaTCu7S0FLaPgVJ/9UTdpwQK/JK6ukDTp11/HzID+hMn5Ag8gXvEfEl3
aBXdy4/rcftL36Khg6ZpD7yytaEFix7LYRUpqz7uzB1Ti6fpb3eAqDHJ7uL+LPSHgXV0khjs9itw
ghbE89SA02mx4W6tmLuz/zCr042IznlpHk50GALwK+dcozQpJ7UvwSsnYDOgg25y54FOjYr8mHQ8
ZDT97ztiFbcguG/WLE9OFhGN07a8MGOopqQte7gqjq8daWBCKaA+wgB14jn45S8EtH6JEoX/WSKS
sEYulfIqN66wdOxEvfO/5W2Fhqe7rL00XLubJSjuzWDsQ/c5peAFEQZLlDydOFpUG1VpaGrUDyqY
WzgO4dXjuf356vuTUHrQ4Y1REuY5X4M2by5nka3SGQXwpve6yZzAoWHnBYMPGTAmCtH5yz1n3PI9
Fg94RT1ONe++W/Qwi1PWsOtYxc4XYv+pi0GNFoyDBzuof4ROHe38rvL7AyrO0pR7NnU9wyB+utLw
Du34pLmOrthtzmHWMgufnv8+lX3r0LBadO6166WArJTEcK7+v48sMlkYH1hcZDYWTNzK9pNJbhB5
Bc2iAyp8Fia+xy7AOzBOx/5LHqvnzgYzx9b35IRBJIJ3o2hedO4HvERSRRhZQeKQxXvpN5JvfsCt
mK4/zWYbldwQ1CBERjBNgqOxTsSPlRuf9Eg3Q//WNCOmP0YtWqEHFK/s2A1n9vVoeTxWNZvKwkKZ
GQnsBikLfH4EQjCpJUD0YNj++FE7qJyOLlFwnIZgwa+K25/VwUuPUQmTYnu6CWw3MWYdfGc9MkQo
XpA7KsE47Cdxtw54uMsTmijw7WRMyrsz2bie1XbzUIAWpDRebSathrcJqWrqwgWzcFJVlG5PEfhR
u1Pz9HGgihwEtwQp/yaxnSgOX3xg6wwg5R2DFLH9k+5jHcCH+roqPXu+9g0UL4UtZpzwJWr71yr5
js4wFEYQPPCC++mqUHfhOQnGHFQ3PAOm/c0TBrRR1b4CwhDphj8qWuLPwmUrrCsMTlJ/0E0+tcVd
9MgORek3gE2i1gJpgI5TnnBqOe0Bh10VcIZNzOLsdKLB8PBW/ZU/aGIQqUpBd8ghGJe3kmK1xCgY
hfSAKf4CieGqJWsU12vdMQmz6uIIVE3RxGvoEWkW0pNolW/W6epEqnSS5Nlf8WvMyABEedfY7tSy
sN/SLfssz/rCgcZM8VLrSOpw64XqnlGsPXY81zQ6XSSJvZI6e9lBygRpRcnOT5GFlMO/M+3v0EGk
DPaumvf0XYse5eg/885qUIc1phglb9Xy0EcrxI29OYbeWoNr6DxNIoQaUKYV1WkVg+hxvLgyvgxH
zQEBVetK6L6PlT9hBN9TDOAvFRyL43yogHQwM2q8fof7n/Z4w3tTA0+xN8LTpzlXD8BQqNbjbTw8
Iw8y6BzHQudFTYqI4lZV28GIhu3Ay5yKBmOZtGkubEvunObuVyYpibVzdJFKatxru4Ukaht/6TbP
V5MYHIfjV77X00nDLWGeHttbdrlQ6jvqfFFGnDK0rMVjkV4Ekw7dY4GGFxX7gAqq9hs1MDlytzV4
+6YQCTTlE0y7cykx2GLNqi0HCTHT8vNKb3SrRIuTrYx3/dMQR/5kWdpmF+14fMxFU/+cSb34z1yK
41KVp+J4UwVy9luRoPGYB/NhykwZLlhhEQdSgcApH4ZE+U0mmfPN2jx/LFH8dKRGF23Ve6fVn/8S
ssqjMZThTn5BZhG+CshuEui6Ra6qYvfOxdIgQ7I03ifx/Wmzogx2zm1peKGw+3AAtQxVovOqmOMG
iVhGKdSl574zO1vforKKZDH+syUdtz++4ZcbTJKDN2E+xfEfIK+ID9qvDNZ9CZO+zUqOfMffLtEU
+UyHnnABLdxTnDa4CGXbevv4pHnBkFBSVGW2cdPtYmPgfYtz26BBijeVqz4r3KJcvMT9FnlfN/Qc
j9fNIiKYd+88y6UlfwhOwcO5Wte0dDchL4J/R/NJCgYdY/Fik45j3/zLsPfP2D0AUvJZ7akVKx8t
uiReVUt+xGoQax+p817u+laTwJpGYLfk8fTePUbV/Sr9vIFWPjLl7NXBSB+SDY39DHb5ygr46dph
3ZLgsMebvdZj9fRwkVyRX2i1xkoZt+TFv+NAOdbsJfQivdk55Kx0Glh70BwF/cE0jwor75KpXTNd
jAfY0n4TMzMtKoqoTu96jzSONy3eLHFsKhXPbqq08zLoMemaxsc38NYgGzm+ETIXEBTu7QubcTqS
5bFxFneoPLAXyou5ArcBz7i17/Cvz66DeTIYULY9z8OKnpsMxapu9aZ57Wp5TuynWng3yiCJL2tz
wvgFl7ReaOtshhh3ylTx1G0IBXv27U2OcbJGZPYdUsZFA+2oiFTyV349AYfsPWTZh2FsksmM9ao1
ooXlxybJDh+ARm+nSk4XgocY0xjGn2iLuxPmtqyqB0nOCnIyqqxOF1FpGn8WHCusjoWLVxpVdGvo
IhS/hI4uM03ZA2inVhtlJI7UhxDf34Ke4nkqrEsMDhqf1tipl1Q5HEDDZtFZ1bpfZh7/w8lPKh4o
2JdY3sGSowW4vn6WBs/1VcFZffW9KN5kC9ZPkrcTAr2G/GbbhmPsxD0yMIXZYKhPcY3QzQEdD9Xq
fsknztSel/+FC5hp5n5U7oOXf2CzCnnxE2Fiy7iLb0rAN/wrpy7c1iDiL/WyVaEQzcch0FrB0OES
vgvAAdFiB9+95oomJVLkL9Goyu25ir7eRyOqowvNiRB72U/0Xq3CQq8uu4vuhUOjv/KhJGkC7pwN
GJAYt4pU+HfGNXgr4+altk4kAV/TLTBYrpCpExsKDeXiEIXZ4uvkxkRFg+H2B97sp49wK7stSejy
8YErygNxW+FBJEV0XEYZAdklXxiJBDV4bL4hLyENHx1RSd2ee+GX1wRVuiUqiyKdTk4QLqFt5nfj
oD6I2SB88vBaJma2Vn2DR/Px1ZA7DGvPynPQNLqk81+1Kmtt0J/CrK3Hcarw5F6dlS8nSmNiBCV1
r+ncZK/DGmnDfSbNGJ41PVz57H4K+SWXHrk/OEEZ1ro3Pa1t3Ichup29gRUrqruUxTF0HS8elKGw
e7J8/Flmwa32vWinPUdVZ5w1yD/9tOl9vUcpiUsn2bWjk+NzCSFqXrMI7u4V+AXlZBfwyQGJi+Zb
mzT+njz9fxjUWl08IIwinQ/6dofTfd+wF2FuW6W24mUzfsgXFyktsFQ4PktkS1WK5V3OEZY4xwuZ
yR3Q8yD6l2BIkdkkxOdm5tan734Z4Vv/7IfozAgFNlAdkxWm+Dh43cklwqjhfmfvZuucTKGNgfrL
Zc3UU85mfJJiIWJ7zAWNxKDsRD1RQLW8+25fkk0yDxNQaloE5D1Hl3UcoFstIyKXFuA3cIj0PdL3
knLwWJN+Yn/pveIFqV+qti0ohr8VGMhx8ZGCAzG53e9dTj5tXvrDu63EfAS5SHOvVQeUB9JNhqQX
PVh/LueD5ENKgz+6AS8HHRZ0Ow4yrxU3Gt5UgEwr0b1t8AaNL/NKjJl0U5nQqavF6FDV/dEH/OwY
MW6B5Z20D8YNHJ/EthqnHG9w8HIOM0bveEnjapaRf/fDRoY0i2szcnOUDGcgCfOS4LaBce592sM+
nWPyLCx99pmNAeelTagL24bHVLAnNNLhf7jG6UcgAGPDvV3AeHsCt6IA/sraMUv1abYXf/jMMOxe
zXSAN09DLmL/yoopAzvgHVstEWWiFu5ari1GqUcBXMN3psfabzQkI1H2K92kd5cIizAk1KfKRswH
o4lAWDH8vC+qt4R8mOinECu24IWHAVPrDfEfGrarvCCMvQVpGvS42A+2NfqIlOYKXmlv4os0ex/Q
8A4VhEqzw8WIU0XJSueHAi6ux3BvU2VJfReXJde67KENSdU7qd1CkNZZUi+7fjgYVaYSD7ZltvLC
ytN4jgBnzJVVImxqxtT9XIdZco6t+9Ch/7NjK5wCrDrUFz9LKtLbPEpzSGn/JernazCmhzCL3+4Q
qSyzvphDCn2Z0qPA/Dsc39rCoUoSYaIocXSO66wW3YxAPMwR2w8xVb3JExdhtwBR+FpGqNKnRjMc
NF/OiduQX0c3LijGVm+EZ/a16/PSB5pNpx85J+9zKAJEkNU+zwlAU8qM04SVFfIV6CigLdmrAkT0
VOXM+maWkbFck+/ba2ROvJLODEWNbTCsC5lwLGvMA8FwNvJEhkZJShjsflw4kSN8xFOH537vy1W7
40vNRewT8G2th4hCfn4Z4PmEdNbQXH6xY34AxwNSEiZxG1uED3Qca4XaT5hCLuzoki4Pb30uvvS8
1uJfqZZ7dufRn/otl1KSD9tsThxRr+ciNEvQNm7VF/FAV4YV1v6LntfQsPgQIV09ScLuoFt4F5KK
eE9oiaakDpsDN24HKEw2mva6bQelYaeKva6kVkLQE0wsTHwpKxvvuYF0UdZsSaKSnVOI480VvSMU
eNkQLDiT4nvwnRcuWojnxNG7WOIBc8RMfth+6vm8MMzN1dNbbVWP6PmdwRuZu4/ehbn8P0fhpiIn
z8sIoyeUR88gU4r4wEBKSS7rew4WRkv313wDX+gXi/kdZ7PHFzRYYA+cojGZFYIkEmflhB4/RMfM
MocJhLkxakJz9oochULWEytesCeIduuBfromhj3ySTZOq3N4sEkk6HG0RbsBZC9abFbsy52aGbPE
+0l1eS19oJPRABsAf/mcV/b3xPAyvziVjOhBAExTmGiZrnM32j+qhaKVEisgps0up3JMRQ25fQUY
kBLtIG7jowQO0Wh0li2/glzqLqFjEH8SUxawAEtLaTjMbiPsTDuM57ErrjEYUNtq/dLwtq2bvGH1
8lN53pOuvXREErmJ0FpQVYRPgc468ZGVRkPj8MNfE1j3RMY1uivoQeUvwHZUREbTfTlOqr+4hgO7
dqBW9IwW8PaSlHNjAy0ZF3BDdYqaMXXE6qmO/6+FnE/d2lpJnxH96Xnn0xOklrV/FFn1co8k7KFc
RgINkTUYKCUmZOihR4Zh09tvCDJgrAlQKrOceQHb20IP8ez5Wf0eupk2I/ewv0IvH2z5fz8iQ+qC
KvFLehUP9toHUAFhb3OVBxb/npysoYxgxAhCCb/03+POJlevjw8KvlJvFxBTVFRAEG0XIrZYcAYZ
LwMw1GdQWFPHrt+ZpfcikL+anqwCpP1zSvkUMQc5R+7MMdE1f/2z+l6MdXzwVyXdT/Z/PQ1YdzuY
EvsRqY2RKX3A6E4zMxm3ZBOP56kph6O0KdNk+RO7ulDCo/abUrDLjyw5xy0u4psrvXc5dCKBwprh
jwjbtblhTKmZjcGtpD3PhP/ahb96bh6BNFmDAWwOUEDXttvDB7E+qO4P2xNicznYBsBmBRd1pDmD
LUOPHsLyJcHH0FWVTSRA0mCzXvPCnfNuELS6VJgSzMcueA7k0ab2ThFzbppBiWnXK5V6g0Chc/GC
Yg7cHawS94+x1LXspKHZWWmpAwDaxvA5htBKYCpczE/viVnd/W4yN1vLIJEKudcEjtFy6VT4IVWv
lJzB8C0XtrZhHljZtzb6QdQCjaymZ1b1BwCmVnzd93QFqFdp1qrF7oZQJloPJltWClLa3l/Xv1LF
5hKwvl7nXK21lKFcNfLK7BCdCF/BJf9SwhtrGnwWoLwie8GnpuMxi1dZY4nW4uXtPYv+SP+gZAQm
5NoRomBqfaAoMYSDlCz7ngqnZVOQuSz0GafuDRGfxo8rlE4BUvbhuFIu/3wtKT33xeyDR1S+Q5Oi
qwNz1PEZM2dvyM+jFPSdZqSFheJNfxzhTmuOzsYTmIVaQGLs4PFmIVdROdjebdJULLFIw1RaBeF8
1aY4Ta2dQyzb8LeQmEYJK420uv3xEWyMaGpR2gtfPGDJO1E+SrP7dZ2hdS5tS+FM227wsIh2IZx0
NLwVkvrNlmNb7lnnm+nxDCvtYxRpjVqoLvcAZBoPXnHo25vUH1UNo6/LjmM/oaE05/erKl1cPQ5O
aOujg4TosyEMmRiHBiMFTWYE9VH1dJlKJiyvcAPO661qquV1p9wF/+g4OnOpmFbP7g/RJD2XCz4n
g/lbFjhDTrcwPM4ykk+wFxwmsGabyFCdo4MJLVo1v1DsWgTT2Z31Kkoeu8/1apXLVz6OdebqwXgU
g60na5Qbx1HAg3w2k/OcpjPCm2LtzxBVxtM35gRBI2k5oHqo2EdlfM4L7/lxzh3wU2+oV0Dx7+dX
DJ+YjuHcSqEKTyvIQWZ0hkmrgYLN/lR9hJw7jInyQ+9LUT5+OQvLWYI/D1Dc+jNniwkxZTOpA4HW
S0zmP5wI7bi9rQvfVSmdweCL4M5AQtI4kfC7VAkPztiZklOxjqqEJdWcf0ThJJcuVp1odqWE9lp2
AE18R7O9JjEV4XGHo/ainm7vY1K9LB8GkZmrtTSbllNLpAbc1MGM4q3YWV2L73zy+P9+L1H7V4Ch
zJL3H9JtPV4b3OlUh8JrF1B2I00vcnjRYVOhc6feLoYqyVraSKj3Fx0nuOia5Em78sg80Cco8vgg
S6kK2+Dqt9Tb/v6yDCeJgC0hyroOFdGPxhx1qml6KJsrRd/7JDr6PvMXeM8QCiEjKoDcOsH00WQl
X9L33jAe4mFX2PhvnQI74+P7sMeCLUrvk9bfb6hkmtWp+VPwmgReMQgPW9CMKziOpmAHOCuMgDfH
yRA4HQZLNOkZtGOkmMG03yUO0WH46qf5vxVStrZQMiITmucyWM3H1ZiOm6rs7rWiIreiN2y/aicy
A5Hcgu5b6xmLTV9GmlcyK9Wgr1aYBEyPr+0DoFiDwroCM8dj2VKKFTP+NXTeuVqKvFOEaT6H7SOn
5l6+rjI0TAcFBJiud+vMDaLmngGoY0H/0FwYY5s2Agt9+dsmzqzUSKmD07OaVO5sHr9jnQfHY6LE
lINqL2PDgnhW7E84jlehF6KW5d+QIFhfAksh5oOjKqOO8mSpOEM7+Z3FGWQiiY1OdGMFBe378DSB
ynLxDAMshGcvKTV2Mh2wgGdFlzXSIiOlsQjQt9Pi5QJnT0t4LMCmM5As4XB1e+aJHesRrIpk2uKQ
rGpT3Z7YZDO+SBRNfr9BgAGGEX6oferMNJr4moCMvMX8vhIgZvDZzrU/Ua41PzpOnAVDvH4Yc3Ek
gbR+ROx/pNMSaPeOECu7e195XD0auQpYp7Pkfol572cxj3M2VbQeevu2BmMdJBP7NDC4CGlY4tcb
XjtHKJiuMhY4mjf7vZd/m4VEGRt74UgKd6vj9LhyAKSjE9yu8IBucGchIOcoiH8xuDAGlhVmNlAx
Gn+0w+apvQAnkh9AfjHGZt/9qduW/kITfxWd9MECOT/laoG9OufUw96WYn/AYcLgMU4wjZ6gwxtu
tQuMAQk80w9pHbt7jeB5AOzZeGn+tdvJC2ZOcqn0ii3eCeCvKM8IkCL6HRdiX3ZP7qFjI8pQFpru
Hku2AWOXO2rT5BlW8QopwSda1rEg826GvpVko23nwRo8SqR0uj1mM5qh3upcNQb0+bQcLOOjJHYB
5suraPpTVr2OO2s/AlqOZ89RL72xe6P3AizKuHzNNOMizeMpMIW4hS2gLz+bYPQUdeqoBFW+tukf
itBkikKTf4hFIE5PZrfo5xxxOPtA5h3tQyDEYQZGTejRIWC4/o03RT9lNiq2SJ0YrnUU2sBgyLrT
1CT1yAl60Qfm4Fic+e3bmcdszOS/PdvkeUc3MTDA1Jvcq0+k0QQH6sZutiW7vYlqPNuYyvSzVp68
72glqawucuoPy3DfxjYuCQI/9Xz1+OLtYG5MkRAqPt/FNMdwGUj6pcOUNQyql3wZWkgVmVI4M74M
gjppuggieqpu57jaJwkRP16QDKwpCENCZafm3EwxaNjKd9iEcKAAmBPjsKMe+/VO85XuocRS26xF
mD87axRqEHbFNAvFjUfMVyoSl1gSx85iyl1e8r0EH4anpLFpCKewpaBC0yiJCQyYbdLMaTT9n93N
lJz1Yr8QbmICsIb2EhnxByomJn1lN0bMoohaFrcTkkfqmjz1AsE8PvloQkMjtLIYWDfY7N6xCG2r
N6rBYhrLipbdx0JYLV7Sp1xI9AmJPPrXCa5FmNeIL6Yt92GSwcdBqIF5NGA+mx2DBjFnUL+lxFOC
9nApeihFv8nJ6XD/i3RQ3bRSkpB0dqGg2rfiGc28TFInn/ns+MVL8Wz7eQXsSsPc5J9BtaKeI7+h
HijSpJ63BFvSYkMgB6XwYykzpYAXTK1H+XMeYJDycjP8QBL16zFZbkobuq9tXu6pmcu/niAA16nG
u1tZq0dpBuJqFhLNWegdXHaLycnLjg5FkNpJmeUIRi6YFavz99e7FLZBYJo0aCkNwZe+NLwQJkKA
0ZkUSgTf+UW1gRoI2T6QepKkcQ3UKYvD+g8alutsvC6Tqnbk4i7K8mYwrZXR1OX6EJtsDL66WdKC
m4ztFCEtqyg+zQmf4vVU1QqIX/H/Yze0pezLB7tm1QgWV8abE47oZkwANnSiu9tu67pNfSMjF/5p
KosFJ/JG2qNCJBDpqjhTSnH1JM0WKG2cQK5E3KD9nQrRH5P17fxl1psShkFUfvRhJQt+UfZPsFCj
vY4J9QVEAL3dDO2vJLthZrgJ5CgK6Jh3QoYRgLw2PNgpER3oYgeQNgIt1k2gJd3K8rm2I5a+SDbe
r8JgZKV/L3I2t9LiwyAqSTSdN2hFK8t8kDaYe1IohO1Fv2iFr4nQSs36hEKD6QyAj7RI5DLu3lRI
n8szMtJjyKHSySgEdXZIudOILGpp8gepdzRzbJpCtgFwsi+s2z5GB5vly7NAEgaBwEf3BZUQOYgr
R+MeYwo2CuMh2z/7qGZwq17rQghpByxiwwrba+zdRldd0zbVeQm+ieLtX/bnTK1ga3rR5Nl3V+GQ
UDBPFisW+ev6deHsKp8aPYeya92l9ooTukjM5NUZHauPSzT/EZRv7Pnq1X1hz6j2vsSO7C/uZmvX
TGUYGNMnD0PShACMfAS1eIrcsI8GVqEtb6d87NTCoX6lMGeNHxTs9XnwtGaIvWAbfDRhg4iPxRLq
SLHU7+aVcdIA1dfHpEIXcYTM32LV5HU3y1LXch4IS+Ic3nSQuDL2b1BtGpiB8E0kKIid/EFUoBo1
uQ+eLFKXFUaywGn2gukYhJo9Km3H3lLtuAWd1zM8iWe1ZbQ1DL3teeHJLkJ2rbIQe0rWplgJSgOq
Cn+KQgpTK0xuZL28SrpfLK73l/koaAkcjtKyMjcZ8ECwqnd1RN7CJvYFmkETaqFp7jRL5A1c+3/l
6JkAj1aKmhYaC0Sf8Me1uf3ruJLS0tCvj88thatGd4UTRj9brfdR57A33XakqVchLLm0wj+7ESLl
bjFvrf8HGwy6vbchXaM8uvwkanBYZMrrDgdrK50X6J7o76244K2F9DFedSGZayv5wSVcAS+Gih84
MQIWW5NrK6PvYTbUB4ORSHGbwIOij8A2/yEWveIGST58EXSwzvtTDID2ZCUQGy6S9B7mKRP+AGC5
hUHTiQlRO4qqlxYxLmn5+gaGvdny6t5Ws3eIff7K46FIWEkVH2fmK2yGjycwFP8eUAenLesghIOf
qkzBlE57lE4nsKHs4/kcYSbFk2O87HSoawgrGMQ2Z8zyqu5TpMEDS1igSX69sUEALAgiifWbthj+
ulvZRjAkUz11J+mrZL5fHjRl/CMGiq4nq+ik+n0NsHJdT7ggep939N/SZUlZZAoowETO1Ca/HrUT
dhIEscFqJc5wT49DCg4u9Gy9Lg40FOFlZjy7TDSgVbaTHk6oeHRJAQTKv22O8SkQYdFsHBZbxQlT
MkLoLfxsSavDnsSo9YMHv6zUQHXM/0orDoH7ZvBBpVQ9zALfU0kKUdsQqnJIksmnZEKvc+tvVoYF
frgP7/Ck5Fn1yT4MZeIbWi7XrYnbILPdkbq5RF25aC8M8w3DHBPh/PjngRoYLvlSz7h4ZTYF92jM
+R4yXReF0SAwGl58xH0pYU0e9Er5c+xBMWegSWnUocDeQDVeUChIJ1C/BReB+0ogsKew+4ulJenT
R1RNjQDkPMHXaFrFbft/C8mKHdWnGfbKK9Kiba8m0nN9IPnkNGrnjUeTzS4COoQTDYbbsuU+lxhq
vd7kwPx2WmpYXEK/ZSV6zE3dNYjOPJerzlyOmpAeLIz6IhI5/w7bjfu5EnB2wx3r7IGsvzZQu9da
OfKjwVa9lIgn/zweloHiVY+z/ywwvZSUED2/7Dvqdv5QmALXwhil5K3z1kzmcNC5IqRZh2zHrQEZ
0/7y1YFoPqpvFwTykhfaT9TjEtOUBWjKBXF3D4O9rl9IwRun93/upNn/u592Pk6PHxXP0uvYdRLy
9EU8H5kPQW+Wk2qTuIv34F22v6CD1tEReZTUch1/aYDjorVd+uaE9/Gu+PT0Z6BoJRNj1pIm+bRT
ewPohSVwbMlJ/CRV8vbAdUzA7Gzqy2hNlSQyzWdVBNWWQAvQV/BNh5tvLja07saWBJ0A0bo0XxhU
HEXuO3s2TEVqbPwI9PPxHJzCyFu5FHmzsZVxk1KOIzs6FzPArq7DfiY9oP/wcDSO5xdEljVI7mov
uUmV3/hEHdkUz7MkABqW1i4sUIc6d51KtUGnjurb0uB3K1vfXgbdlx7FOr8Gno6Gi6Bf3j97J+0w
ta67yGXp79Gp5fIXbieo7FuSqFivV5apu27QIOHPzeiirmM4GTPBP14wCxgaxcW3X53KM/BSqUHr
SRaGIcICeT15SsU/TmoOwxvHMlM6HUCfoVF2Xlk8AVnyhE7xZWWXY5nzb+esKLF0l9wqsLdj9Kji
+nMsLnWtDImudCQwBnvekTPQoWfIcLdFZScWZUOoQVq7rc/N9QcMyeLLkE7oZhe0qk4t168cTyXA
eHB/AZvU9noyddMlJn3R9ICfZmirotPg4njDQm9J0gtz3fB4HDKv30urvkwycSe/RDpxd9osnfpJ
x/+UmSud0YLn468ZNDpHxkTTTC8tpTeDsLP2mEMQF7HzkqsgumLQD05cJP/r7/tQvxNKhvIn51Zj
xqWCwyEeWMM9sQoaLO/ioKeAgDfOLjQ3iiKm+LVfJnL87FD2uT+x7WlwisgqXPH8RiD2d7l+jq4e
xe3JEh39x9DzCA6o4kAsEeySJKSjwyIfCcudda8Sg8+UY3tf50z+V4bJ+0PX5tSpKLGOx8kbIvxF
y5i+0gDe5KIsM7pvHqp+9Wp5J+XUEE+Fp/JKWm2jYRjrus5/AA/PvOf1hY1rrzjTip+Hi13zIdGf
NTEuFLUBvqNmq/Pjr77Edpf+B+ipzcqmbQbUq7hv21X1Msjv6D0yG1xI+CPLQDgWgMuyhQWVKoT1
jKkzV9vJCnbF+EOo5TC0WZUBvzroR1kdqhcZiKdprzrjSFDecbasZxQUkTPssMFqk/mQqOw5dUEV
gC2rCGsjPj3wG1f6CadtJRq7pQUMjVP9Iob3MCPF8nbX1mWxMmBQYx1SDlD/S3xrPBUmrXiN6FhG
RKx6PDIY/DI9l20UwfI5FkZbTSkpolayCNBooEBaYMacHIEg/rVQ32qg85CkNwAN+tLEpoHBZMPe
t+EZZ8m0VSa6UOIhX0AFuH6eN1riLzci96iX57gGM6U2Mett7v0VJuF2Hd2YpV42W7VD9chOURDp
nQUtzasCjiZx4CXSCIl19uJZrnrIZ7UX9nHBV3c6qOs+Nsca2ET1bovocpwovS/0j4Y+TiLkDK0a
0PjrhBFUIOKHcFShztNLEf2J48TxmfqKlRRDfM3bRKqllf2WcbPColGFqFdKqmJyBCh9Dx6l4QLK
kLZpQc+9mpSO600v7AvJp9n2/L3m6fA5cwGXsh+WksMbV4m+WY2CCc04hUzZibw1kt7pUhVQkSVN
BPh88xNaXVmwp4oPzEsWakOpZ3BzbwF+c/3tdrIzhaqmEDWpkn4dszZAiaVLw+mtoaIPUOwMy4gq
nagcB8J413h2NWCRtEwwvyUgBWUZZ2QikXzYGJ9Tga3jx9T0Iik4kh83CoXnrJpIiRI+E+YR/nsF
8RRMd5LNC+llnRqKVsPScGmVnb1GijWzwBe30dZ6egRxFRUz2uAQLsIid99tzsU8LPNyPe80ZN00
Sz2H1LY62c+vG2GJxIFiuwvur78xoGqPP8JqJQW0Htp8gtJmy+aggNAo8b9bgyv7yO6tS8VQV2ZA
glDBU/1l9zf5e8SSgJjiP93AZCMm/fdaucJBZORhgGXkFMQuJQiDG7gNk6N5aWQQpr5kRXeQtLSY
s2q/vjBF5K8+Qg9YuQFDpYBjw7tuOwlcnLCZ7dFxogSCAg9mXcezA1HD5aLrVb74ua+r+bFNYm2n
1NOo6TVDQkJ1kCm94GbaC63jFQXGQ23pouaJedxb2H+VcILkwKP7F3/0VPYfY0/9wL2RIjsVBqbD
wlNNIkd/Uw7J1xhAxwGvxyp4SrMCxcqrYPo3xGzOKVeSXjCDwj1qK/1VSHyKfj14N0ExrVaBKsWS
X00EnL0MKezfzsHvRfDN+co5fBjM8UV8FFzmqyi54hLzy3dp5bKfvsiHYAsO1BfjAOQlSNXJ60tF
Ipkz1Y8iqjqkMzasz84xzTavMzUNlO/ML/CXKa1cy0J9h0YlN5yw8vW0BUAJeqMVcRs5X1B8hhsp
4plg2gF/g3Q8C3TYpC1UnuFsi+F4Da2gfB6CciRuRr1WikdiJaBplX0Vs3jssAWDIBxucG6emDIJ
fpOqxwBbTu3PMsjPYKixzKcqJ3wu0Woh1QT9UgKX1nNw/tN9og8i7EgP00XBl4ZdXeuWqkYg+2+x
8aErlxwYNLNdtCDZl2Zs5WBOQdnaR8OgjdF+60N4P1+SdQ6thjSwR3rXN4fZ82haczrZerM6zlkw
Rc9vIazpLBtgeII2byAqnaDIzgOj7TTp6H8Dc6EXjufEcusdjWna82m6I62GiPb5XIK6XRHKVzmb
C8HHG9b+kvuwlchDD1m5E/YM0bULyGIG1jKl8xWWd3DmnX4wsuV5NB6wbr5iXFKiS4MRck14QUBa
QYjzLC6RacslXhZkJ4nCNzOfn+etpX5h2iCEblf1kO+trAowIDy6uQTam8UwUNgzPmIhLlWO6M3D
ymnY4Bm9wv+uxQQzWTAJLEGHrwUt3DD8nwP6xaJf9NYo10yWpLc+RsawQSns0HLa6249YF2p1QIy
oJ2bLum9uTIq+LaZ8+MYXj/ielYhm7xLyZB8FTEsxhY6jryzR9xGgBbln/3qcZ5zytPsHd3snBut
+MVTMFiuz2Cd3bpb4BnonVImu6wXf+YSVRROuDQTJWvRobOBsBe1RGVZEbfdl96UNFDWN/zKTmwA
/xS+QAaoKGEVcTlbQsn1lbc62ZLKS3jkUpm1xbS0GsCuplWVX4H6WPG/fJPcWYpVAyR5gvLUSp3E
42Aoj4xYnDC1AVmiC9Y9LXOM70+nn5G8YclSn6qJii/KW8aqXoucgpX2fuvnqkba2abLu5+M6alX
BkdxAzXzBW7nfYLkfAgoKvCNnD6WVs1LKiX/K0aAwx/Ys02XolhtFBwcvBr1V6mIKHdOKoGG0AHz
Vzvdc0yqFLOYy7kWWnYOpU9glYUV8f2zBTtlBzNpWK0zd+AmBLGQSzETt24BL62dUQ79zvJj/ibm
Pu8bAUNVgB5t8JHTTQQCoSeHdQZupmZDSjkZfpsJcCY8ek0h995osJz38tkOJM/oI3n8ynBTDEe4
eYF7w6yYM/jugVeszGWJLON2Whe5GZP7Z6gSn2z0MkRKo2D1qztF62scTS+9x4zovbLE9NzdK8sz
tkyTsYjB4d+vZB2wRsmgcI6vuBINOmhqSCa8iGEs165YIRHh5MOcdkSG78J4qlKiB60GG/8ipvuD
rLETJTj5XsS8ubdAdlR28VlIX9O29NOWfpYXT7sufmK8pCQOZZzU7vACn6ZYrvBOgGe26ZA53NCP
M0NsFVAb1tcwzINxCcTk5dIcu6fPXjFdYIiOmAKk6vP38xyCqcGeOb+Ck0VgjNcM0WwCHZM99Pa6
l/sYJ5rdS9zrAWenV0EtpGw0B8z+yv7n3u/mhxNpEkThP73mWGooffVh6+sHQm/hxBPn92QlbVWk
0HvL17GvLKhZY0TQ5sF7JjtXtbM0qDG5niuBDbKEf4zC0iSJif7Rft6g4LTABOHJD5KVbhLSEHqH
dttdWcoame3DfBzU2MSFHk6EusqOMTuWUGiBUcmP9tboemhGV+0HQKPtTFSwfy+8/+rJqhg0u70J
wdgFvTzLC2v0baHENsRFOjEPFZ32TWUHZu1W2vlhakWZ+ufOm08a+az04jUT2WSdBSsSen2rxtGF
is6HnlG3vljOspVMKCbiFoUj2uNbIOEl/iX9s+FFeeUwD7lwwMQxYm105esHfgMxd1C6vdatm32S
MpNqc4UF5BE5m1GXebM5OPT2atisQpfKI+H9VbXIH1KG+GLTk0zFFCDwrqr7UCC8ORmtGOQEaZ4Y
cRUkQNmCbzZw3OA/fpfAVK1cHE3pg61aSR63rp+7vUfRiKLEDTbU+aievFClWn4zG73TL2gH6ZR3
KlDKbWIKVDAtq6RlGr00cpQKGN8Jb9eVv7zd7IMk+tVY+KW9aR0Ppv0Skx8YQVK+AR1f2BHPC10i
98dCfYetfEDUwFkHDJoWJxdlaIJ6zG/ZTh5OG0jmVEOS+fKYWoXFQxEO4KOLhNmatVwStpbp2xZQ
YBV5ZMzEk0fLJBhbr8XphI09sEvvvRwiNABi3ZP2KstqYuW5f0mJVzkEOsX5AuX5QHCVdNUIGqWt
JEYrnTmDoSQmyfwKfccV/XmFj6j2sFfNKmRjYSjb+rgyZ/0ba+R8ZYBorKhDk1eZX3UAvi3DtwQM
wMY/bO9nHydvCig33LJMHmQchGM4IEEZznnPCanm5hcS33vLnR49buDuSjLVaQy2Hz6DvUOuq2QE
W9ZW+khGS2d+NTVpBIP9N5Sndqdndz8bUPScUs1bZFFj8wQRvqyUERGWIw5ZKXY5xZVbup0n/P0q
ujt/YWzhVom223gb5/zcUMifDIh9JluYuEukp3Wt2r1Y+0UCQ5Ux5N3qsY6NS0hUuZ6kvTE/Yf5E
aF8EyG7Fae1NYAgu9fkcrlrkcXW9LAzdoOE/ZOHYw2ZYkcXPwyOug4gBZo35rawCpdjAOVz2coo1
AbmyAqmvDh68SO2aVhPpMS6T71IYfsS1LZ4anV8acTWnnBFDDGH3mjUYofdCThYkqdmQCSw3vZkp
qEM4e+VpD3mf/zMQqgmCpfjkbg9tJeRafzoGyl3oA7+RH+mZxM0xlTn9HlBa7oqW+eXp1aC0iABG
4IJu9g7lEA8MAymRO6C7zvTPrm4/ixOD4KzSP18hYCfzE5eVPqT2JtzUOWSZFJIVQU0K1g1+X0R/
X/ZQRmdUp0oSsySCakSJkK1L5rF8f12sPQAnsxT6voLGy4PhkeuDhL2ApwUKQPpBSjc94OJn2D3N
dfP85IqaVlA0Uv6OgCwW9y1dhwoDy+T15Sg/ISaAZANsWXZYPTOUsvy6MRwv0gCMZOabusIgsfT2
5d3updV0TQj/yrC21Rgbr6+aLxzy87iTf8/KUJvqbcFi32mrU0LihOMtMYYJN5LjN4owrKg77/kS
Ru72clu6VfoqLp+i0xzU//emJ57ncwH2Tu6k1uI++jDnJ2hBqzZDNfQ5bVtCG0z09jKEw7LP4u8q
jyxEaFSiAq+cd+jOUHhmTE1RQKoG1B5Lxvs61Bg0460ODhnkTHfoihjbZrnh4/oSFuoZJlFs6WYV
qUCWQYUuDW0/9XTUrpFot907zYs1jbeRgLkMlMTgXEYTam/dD+QycuPpv8BKsOfFD+Ns0wSamBHG
hMHiSrcRVDN9b/XjUTDd8152hYfhK2I0jUZXPO3ajzUbJqFTUoiSQRxdjiTYBgJMjyX15QXQvLbW
QHoAaSQuh69I6FOJCMg9fjeziVn5NB1h4+9jU/vL+9UmWYxZGbAun/cOKCsCiJf+G03B2OzzvZVF
aGPJ6+CXexNJRKpyGQTbf832Ymwt9c1US/KwzY9yEervq7wc4IYR1kbUZxt9bTVhdtpUbBBpQXJu
qTqnnCyUIjbT9i0MbeFB+6YZGmg4FODhSoja8k+0+XpeiHo7Dxy9zkkYNky+uOLIq2w7W83CVqAZ
P6jEIg3CPMHZsT700P8XifquU/aH6ef65YWt8u728DO+Nrn5r454P9gw7/7YLrBzskvVWN69E2mR
CDGT3QHZUk2DJVDaT6cllddh+/CZInJ9ItD6xGiCnUmMD7ck5pcz+AjGCFJVLIL5Xi/aDtAv9luq
8HGVI52OlOcSJdL1Y+E0b1zr1ldJIXCYXWaL07Y6oo8WfngFbiGqWnFN5bvmLtlfVOeJiyftFUwZ
6INAauevIRu0dGC3kzPt/ePcCDEZBnDQwPUQ7dRaViuyimZysFaP4b5pyGwNdR/AxYS6CduT5hZ6
QK+dkprzfz6A2M/mRQCS9drQ0WQWNoAEo/YRfXUkDyxd612X8+SfbZTU0MXk98BxXszsUiMH5Vyj
Gye0LYish5ZLU/k5A/oRezOZ5XoRRjIstTugz3JR4eoJte37Hf6cxjbd4JQxH1FBdNj4eG5PWd7t
cLK4h2eCe6ECkNnBO0X9cQ6+HwokshCEM50wU7dh6mQDwHhLD57OlDMEb6YUAlk4YOtPxmAMJciw
bjEDx+eBcz/Gl3+VmkPNvEOmcPKmaegWb8VBbKOwugpcJRR4JvEJrBT1RqgE92zAQ1g7jNcHUuk/
IteLUYwqIRxXhx1zlAv6/Sfk9oq+WIUyqvoBOpbv9JsdyZTnGaK5JMjNVRSpx0ulm5bq1LsjKgtJ
CesWZmXQSF4ZvGbS86YOUmcahZ6IQ0jvJt3fd9sDPQolpBmVc8LsYAhunBNQB83MAvEbpfZs+1Re
R/7tQK+piMJvb5Piidnqjt+fGV7ibVbCE8Y1QFXdt4eyuEmiJKt9rhOd++4vuZf0ekSmkafkSq/o
8hCKRiRj/lTeLG4ptvr9PDOg1ZqAdN0wzjd/noWwYvhY2cVzW8bSY3GtKkxQj90iu+eAy9PKADY/
1rdGsHWVZViY06mZ2F2FydVu9AMwS38txOyuwyDO/xrnZGAeV1Gxr7rjiMT4h19ZCvcnDzDoi2MO
dQCxYiV2MXf4FHXuTs0UZIGBuqUvIJ4/eZdbIxiSrL6SZjF48pXrcYoQLyhD1SNST6OHHx2sutmk
3QlU7NM7yQ34c+6XjkAlsvNRqY4I6fZzacqbytaaD3AluIUvqUJzynBB+d9dk+prW/VWp1MSlKDF
Z56em/Bjz9H7EpSsktQOJxQfXqxFvBjDe+YKGrphlJVKbe08FwcrUOrbisBtewI6Pt0Gu8iljaU9
nH6cIskW5OKN4KWvU2adyxjaMNvYmel+N5Ey3ZvqCreuoSZEBw1bWnsZCc5wAGrMvPrjyVjgBojc
xOyPeypfkJcXPY/crlTOY77Vdp8jpesX0VPcmk0r6R4liBSK2JykUC58iHka6DuMJqaR2yhnV2Ye
n6w+ClZHmtpBUYQCU0+h4+HQtW3Uk3c92t3MiQhDVc64M36mYTyyKVXDTyIXJ7FFElrovShcofrM
Vj04t+ZQAhdxwA+V6bLh9mKbgNP4IihGuJBGEI7L8cvCJvqGNh4ZvzkeKJDEhQCGVEkh6l150v/B
KcjAd0iLrpA+b8s7oLrV4QNOUjuuP3iEgI7SWK3ZAayB0nm1B0D/nT52WqdQG9K10QOjKJvuBmbG
jDfrjcFZZPGJucayxjfjbh9vZCecm36M+TN6S5bliB1vnECYCap/S2W1Fu0MzI77Smsq1xkyeS8O
vMLFM/3ymoQGLaE6uNTgfBJEdm3pc5yyiryHs6ssFRj3Y0jcRpezNghba+S+yNQ+LsO8xeCzc5SS
9/RPv4ffksxFrCc3eFqMm9A+89WrsCPwnho/eIw28qXA6w8LM+chJGyrSwp3RdAI0FPQEBOuB6jf
jJc99P9woeZvIQSvG44ypv6Nvu5SWWRbUV01MRtLHskI1XxdWvImd/FIrlmhcDzjg6VxiyDufoCh
TbL+SAMPT7GM203oRyHK43AcManrp0fug6WFXS+G8V3MAG8qu0hqxRKFcj8JvZTA/8tzV0AOjRU0
k2jZ5nqhsSMWRwcI2S3i+Z9NIROYVogEN6szRz12/O1zMzhY8OT21ktFE7swrlBlDpuXyr+ow6GR
pcOTjBTHsq37T4EfS5uw2d0BGWIV0hW1+lwFqrpa1PBJ8JQZG1TtjD+q2GTa17nEsc2SWqcZteWS
bdTxAv54pZ8r8GoJILYPz/jhEI4stjIKbDSFKC3HRMMe6pauROgCkHH+sH/72sFVdLGWolwSnIUB
KtVHGvJxfAYPki7PSq8rYzqwvenFAE8cX3Z2kq1TmjqCNhciBjjoU59feKx/KkowF20iV/aMfItn
yJXtdOABeqISXwnOgMwomGgSWYNL1ssQiZ6ri+4vSYpqVpoGMNk4ctT0yab8UyXksubo97vQZzbY
L8Wkjr/U5iI/dOEsHlrbanXvlIPkCQiY5TTD07FODtPvS1mJgfx56Kgc7ky8ZWyELF3Jlb304efj
LrVMAo4n+AhFXd+5oG38nwyk9E7hFtD/PKu8xfNRVsh0JBveGFQOrGL9Fe6sK+40j2odrdztfABR
wuHjMpw2Kj/G0MBR9xwD4OXES/3ytGeEKWiF6ujVo43dFItE8KrGlJ0LMbtmqjiLoSqUxLV0TQcb
brOJwd6mE/4ZJ76HfFT0+1V0xv43o/n0ERLK0QHIhVtDY3++br0tbRom8VZKLpabZsCzQzE+3Ar/
gHGNZsw+aOaCwaSpDNeUtsc99+1J6HJyO5IDF1w50vkfHR3AIDcMwWa8RUcoUTYPH9uf7iVXilJ9
tM/SzdOsNL0YMZwaoL2ZVONMuZGUViMFsFDaBZqXkSMwMzdpUtF930blFznNmdvvhtwodhF3E1V7
hpcf/qvgjF3+7squCBFO9yjuEozad+74XDeEU/Nu8CW83xkjk+7wbMQ5v565GO3kXoLDZpIWbE4S
zbOVyDe6q6XhEhpvrTs29SiEh/aqA9JgJsE2/nNpCdxNNkdMXHAlbiyoUWd6XorHY8x/Gczs5avW
1AwcDlrknd46f7BoF8e3q1IJhRdiCXNfh0H06Cj6yEGD9wAr+RqzFdrV8bWL3zo2fydxtfsg7Tg5
sKq+kNE81OYx8GgaeLrX/POjlXr4/m41Z0XX7Unw9/m40X0kJFvJl5Y2c4ASvDV6TWlfcUZQPA2h
m3mZMQJKcx0OreqKRYxq1vBWpC3YkuyvpootVIZZIBHRGwkR1AceeSnbiUXVQq+4KldoCsmv/Zgl
c4wmyDGr8WR8633K2zuL0rhLZIU5xwSDVwc+wqhLV4zCam05efNWtvhzT6ZUW7kvHuSfXwppt2Qx
gjiv7up9TP+Ohq2E5eEYFzyEv26GFJx01huLaFus8L27zo+YzP4aImBPiSIYDI787NDkE+KubyoX
T0Wj8zz8t+47wZ6xLXa727DBk3fLbTxCXr7CiPDCgjF79QNQHgEoxk6k5pVGn46q4coxUNmrDCjU
S6QZe/sDOsHRSk537qJNdB2+88wAWaAQsciptOgkXDGfNwAuWV2khDPHscikR9PniC+yOsV9MZqh
6a41h4UCo1HGNbc4ipHqK3J4uOvxVVlC+KPhgn0YTuBV42ZMxriJJLxJ+1zWRwmpr3r6ltUvvP6F
bO7YWbMsPn251mJlMjXHxsDeMj6yszlZFshaedvloKUJyqGPSmNxFB7PNh3SYoEbdb921DK7YK3p
aOsGYZ9se7U97s42f2Q50olDLlISBh90CWd3NCoaBQztq2G9A6grHpR8O/FMUrN148du4w/penuT
UPwO4G6U4u9iAPnyU/UPkTLdPm5ESClgOWF8xiyqkPgAFr1hqGvqN7cQXQ5L98TQ3K/3BJ89ADht
hXRqMQRdhLNPMYUx1uhxXoxkyXjmlu8X9x0ETN61k8Yf7uz2O4hrvE4OB0mO7RVo5RixmvlAb96z
H8qfVfB/vzc5gR4IAujpoFCRjRSnPmQTB8UWPDgv4RmETQ6IikNv5K22H2K+MhcNODnE377dkosB
dWlBlbsIgldHuYIALfvcT7atp22dmghHHLN1cI4Cnnx6frC/xLjHy0MaBeC+CMDu5ZlMgjk4nYbi
l2e6TFGahVbtGrHctfvpr984TPTU3nsTcYZ/YHiftqrJ544VRXqGoTcfXc81OWLE+Zxlcla/+Yl4
YRPWwxYTOgE3CQhj0bHeagBunYYzxUUuCYGzcCm4iu4LI3IUXbJMrJDaww3G9ufzCZfekzvehZbE
9CRI2HVp4jMRfIOhhrkbclnPl42BmQmuUqxlj8mctFDQBKjtrOg/8WWzFxXYT9Qlm66o3jlSAEvI
PEWL5fbIyQbzQMDk4qmqATBAYrxtM1l33Ke3QFE6AarZe5CNYintwbfL9exx/MRU8Dh01J9Awjjp
KVDzRV6OPYgJf9iWNgom3Qo78gRMV7/MtvgQbwN/ZIc5N172+GXH1P3sZz6sxqvXVTgRnlD8lA7F
xxo9hAa48B0GgmK9Vs2s9OFJbB/NMjJZgcMJuyhp8cUBggOkIUzZ0lybsrR9mzYzeX8DqE4eqKkH
injBeNnuLhbGCouFsWYSELn0DTneg0gJTwoESIbjU/YSsHk+teCNpTdIigx6fobuSj0gPW/vsKfm
/sLCUz9dSgUJjkgqplG22r+IbIkWspfLD22IcW1GuoQfRizZt58qMtHRPIQz99iulPILpb+S3OT+
lQc/dHsaeOZedBuk0fQJ3pu9LQ/m2AmMs9S8hOhtCtTPDs8eh96LQc1BchstN0I05sWhvNs9lUrs
7BWi22nhBDlOqA6mTkCA/BshAP+Rvm/5jASJCQp5x1HPf/KcRCGjt4rDlvSmfR3TyVIvSYf3Qnnp
QedhMvqPyrPg5IELya9ol6M6WentMFTg9exQbuo822Lv7pdR7APi+oBQE7WelHY/x3QIRFfuzFy6
41yDuWowP8c1IIjsYEjT/XV+wjb5NBTXhxkJ213f5UgxSuNP7CBQSuBrEhbnNSlN72g1r56MKVD2
ARM9V5fWgiwlu8siqs2/UCE8X278jWQQGz6GELqGJtxfgu0JpptTpSAlLbV8+IutxG9dO/Qkwfy6
fu0NgTTP9hsMfT4AYZbU8vjwSnfnWRenEBbg9J5alXx8TVpJYFFSN3A00A6wzneu9aYHSJTE7lQt
SqokBirvkKVgzM9euiYmm9fbiPgxHHsv5/7d3nLHXbB/LE9WCvlyIjhDH+Yb02GDZ09ltGch6Qa8
FeHn5a1fJeDoLbXPrt41CtWDh0AB14a1ZRanaVfNw5/jrZ+00Kmaro/61VhRguvXkfeX3SNpB8HP
R1uwH6A5JOyzlGTmP0/LmcF+dkqrNJzFnH20jPLkeFzed5za7ibxU1++QOB0nl06vJy9pdsDETt4
SKwnAlJVij5Sfb18S1eFvdTFue8LVFIWkz6QoHFUOB4sB1g/vnouLuWSVMjzpzFJmUwKjUz9hjpd
ZI8DZF19dq+gFj5APgPXZCqTjE8FEYjTSqj4KbHJSwP+Uo8a+5nYZBd7523MmviFuSi4RDclfX2l
/DoXsQ9hOUhIhLJHEvQMnChi2YaJ1z5ASo5ViiVgri2JYND95Jb4QaTV5rTo94cB81Xqdyz12N0Z
hpAPU/hPEp3T3N7OoXqJkwxmrOq9pMNo/chQXhGmhVa0fSiBx4lg38CPbnQy0uazeDfw3SveQt8d
1/ZXyCFLn3g3UnpLDlHPCgLYNeTVD/oAzUWh/8scic6xJEfYqxSB77FOOR0VCGuFxqncolzCFUmA
u4k1fSLRNvpxPSamPqLE7rwktf1SZszx+x2obpxAUCJ5ZlEKCptLaxvIMocydZevwzvEr+Vgnnry
HJtaxdYCFJpHAAGEEzQIr+OWHBLUZy1RXeEuwB60tHLBMgEthBwRuEZjp9MZAcLO1agR6PDbu7hB
1kkADWcm4StiqkheTVIeTEKdsdlSkEPoiy0RoDcOYR851T5EkiK/Nwgd6h3m5Z11KDibGbNkiklY
ioKqDFJJJnYkxq4MQIAcGbmbjWOvhkQSkAEMVCx+qb4xuHXfoE1INV0HyB0u1vfZOMzjL2rdV/Ya
MtO+jN72oJ/AGjEXfOy4W4lL9nto88q+2BTZa/t6Yg1H0YJhwZShUAo1wtNdc/VmmyAcuNouYHNW
ZzoRwwkztOY/TKF8If+Cu5D6/1bkpSeFWguNQ6lQDVkgt9i4OByb14g5kU2JbeEihPPEoxm26twG
//kgVlOqUBeSGA6CAigAZ5E1aClqIexblnGFA9ig18E+Qv6cbNcaoOkWi6HLoZSDvQATfUO+Kofs
fO8Kdu+rXTk1kSUygd1xgqSdWL4Fxu48dtv19qTJwK6cSLfha0xzSa18DNiOsHn8f299I9udK6kc
8Gn7o8qU91gyK2BiXwtDZ7ZPb1Sk9R5ZmJfb7uJqrFsRO6NgnQn8/8bAOHEhoDFzHSqBPXFokJSJ
hnXTaNcdNAR3HU8yZghDzPZ65MFh9cRJyVVd7XA0zgMGDJyklpkQgqq7QNfb3jKcuNL5xmxuTFEF
XqSCDk7tQl/OFrFmhBTRYy6HWWXBGPsDaWjInxqEfuZjI2X0w4RR48Iy0RtXmH3UMd4BLEVIqwjs
H0YTUlauiQFlueTLPjD5MYrR48oCVEcjrN1GdQ9dZ1V8CBORtXjHpVQEkh8iyPC0E0tBwMB7nzRy
tLOFAkHMpAr1fswoYIOCBS+4fjBBxqPIfFkHTTorzSmz9PXnqBXQhtJYvMChI+khwgeU/Brj8NeS
GXWD8mF+KKTUyGV/25j1KD0qlRNbj+SfIRaIdm5CFjmbsF5cPnMrFA3E5oxD5vMsrgPTXG08QBh7
QjdjbgRnuLvRSCytoVEiUGwr4H8o2A7+WWdj6KqP8oNZP7XbiwtqxUnCuGpMlb5nIkXdL44EBbI3
/txOLyaJ2rdDOBsbsC4gyX3eaS08C9yrvHIjCANUI83nW4ryXuYBf1v1Y6lNCR0QzkGSUAc6hQ/8
ZPg5BjMDFof3UhWoc3bghNWO83o9qeI03wTg7O8v+lZQOeJtY5tTk/Y+fGUMJ4WpyzNDQAbk3t88
/0Mnur6yGQArPvWJlwtwal0+/ghRisecfXEkAwktRgJ/W0mAt4SCDxJNrofP73h5xGyk1CXHJsfb
rkrFDrRgVnNIpjDJCFNI8J2xuH60+Cy4P1aKph9h8ObFAMSMlHuiYtwwhgHXxCs0oPMp+8+pnA6S
KhiSAAQ8YzPG0+Rjp0mIESximA3qEPQifihKsjQY2lDvD0pPoHnWvcgtiFdKCQ65sChJ/YgjL1N5
tN7IE62e66udGQPAzEcL5tqSx2TK1hxErJ32Y6OATxGeperNTlTqG09xNDyNnyHGYZIsv1rNcsRO
2lXvAmUYPe3GhF/8YjGAcHkEuc9mv6GIp5p8gllVrJ3zMLRmEptA58QFKQAnvwubtEWXi8ubijtY
ADr32fw7Y7GHDCYBJFnjgqNudJcwpZKZimbYlFF6y7C73WPG6KWhNIo7sYMFt5/d4ZmltRHVcDV5
TKSH6scq64plMbp4mptc9k267fI0xQSbnPgNgwUZ2XxB0+yRvuaDxhc5coBH7wN1JDdnI9KqX8I6
RZylsXYgQiPqD+tW60f5kUfggasP94tv0axKlkZfHVP7NNpKkSAzAGbQ0jjB5BOppRQiIAcbpyOe
mB58Fm898ILU0RVXi1kWj0O1LdlVyXXoJ25lOVgkcPupFBj3+K7jq6A6tfVs4aGBrInYOJ6zWmCl
gRl/MqyfswiG5MfqAK0YVtVqQQM4SfmXK+AZQSAPMaQmc6Z9dg5g7i5h9XMCILUbJRF7rXg0MMoi
Ovx08j2ORJ41Roe63RSjq2k/s4/m2ysYvm4c41UHomqHPyq9dUgs+yS0qQH188h7r+OkgAvpDfHK
KF1MslXBNPO85wsBHeBeUKqf7tEG+oipx2yBQ2EjKuZAhrHfY75g2xllYv7/G0YkCENsHgK3fn6X
ETyC9RWcTTt/ubP6c7x2GhIxPPmHazd9e+QBQw/djjkgohhpRmYZR63X7X9PC8S/RT0a+Qw3eyji
k91MQxzib+I8Sx5NAgaN9F0/v3QqkYEgUg2t5PAf+tKCD3xFs/PkWe0dIPdtnuEwHjBe6g2Q8wY0
hvXdufSOnfy+/MYJ3f5RPLm1zMjutr2iqROZDhkip+O8iFW4AUtOO/6pNTzDW/fRiwxJH+qKJr6n
M4PRm+FdS861z8va2/qh6HTWhFzc5HTigCtqVljQ4dnz6yIhtHdoWcvRPOHYC0DPTYHBgpGlbvlF
7eqKBfgTEIPsV3fV1J4tP//uCmBuPVjT+DS7qBAUD2O+q1ZpO/cpMP37zJoNcaFUig6Ltc7O1gN4
FGHZRK6atLQMvdJdJ6hT2HNirARIv/9pIc6vVG7eqDQC3319lgCr4Pp3auEe7QSmV9Jyb4gcTkCN
T2DumdCuucrf2+9DIaT/BhLCBlH6W+XUTBugdVkgkAwAX5ivxiUvYtj3XGWVLsbn8L+BsUAj7inF
FL8hF9J4TGYjvzWIqKKz3VSyEzi6tzG0vT7MfzM7phK5b5b8Yy4hwySKX3kGqAoZDJmpuvdk80Ze
WDNvaMndJa55TCypJucQy02Bfrk/CjEN6hG407Ayn5AkA73iiGUWvZQMTBayb2uyz9BuhSwt708B
r+4MN1TKmFDDKM4Y2Pxk8pXMBRmVUEUqUFCJJN19/cnCZnzxXW5DBGJx+qsnqktA3t07cVVrC784
5/tRpIX49Bv3k3g1slSLec/7dZonqnRgD0VxW2Hiia8wA60REZVV17yD1YZNTdIvuwluGhI6B8m8
7QUX5XbxMUcGhIJ5urCgIkNp2Tpbm0zJaPtTfd8n4oatTGBanWt/2Iz2fLAaWTNqBFbGwdGTdG3V
BDD458ZW6nzez3JzoaGTOidChDXQ0Vc53RuwmIFvm7qdPv4hiiETDVuD3cWF3vWrjAnU8XI5fgtb
mNKJasdEiZ+HPoTJBymJYVmemaR+r4N1LYs905ki57aEsuF8AMAFS9bSLndh0uowwImF0EyycCGi
kAZlDtSmAynKtKxKSC5mcoBb/eyYmcbHsG3AQ6ofYcV8nIss5bxATXq7E+X6QascU6FWfjBDzpP6
o/3WgwCek62KGBixkXmt9qan34AiOdpz4f3iN2JvJ2h3BcU8Kf2Tpk5Z7TEHNaxRi9th6JeROOW0
ecKTJPRxt446vy1Wsoxm74L++SKAMJ8inFUjlEckRwyWhuYkMisVTEEZ7hNUlKMNP/vCNKWR7OxH
a+glwwvmLcMjwt8BYVbKKQp35XhZu8wgDRLTZgdMbnXx3xy6vkZDbpqHGU1lggLV11vpmI5X/Sue
gMmtRGsEKA3lssqBLnuhVaEXjgEzodVLK0KWQMUbJLH5xnmIR6I5gZDFR0QrCtyTaRgqy8vvEcZw
zTi7RLnIBL+JW8ef1ryX5sqwresm8ZVW6yfwepzDve/ARv9NGaDw3m8AAc1z3RFUsXUIpSvbEne5
GOd8XoMWjojquqZr9e5AgblNvUanC3HvxnrPWXJkzGuaYNi2Dq2EFP/hIRnAW4im0OtHpaTSCCAB
2VNoU8Qdlnn9pdFzNDu8V8FBUHjNxjHf/17EmoZ2k8u4cfZJRc6F4beaICvxhmAQAGXgZD1v8F9M
nFWAk7NWziUegigrL1R66xdZhszZh1C0mRWIVZFSDNeExhnvRK+SPAeTZvXzYp7z071gpv23Floq
G4+sAKdsgDtivxCs5lfVy4JWk3qxVllPu/gZOdANY2h3tWhyPW21U1R+hsFLsXkKBlRYkVVbN7ZY
QEoSuFsroBCvY8NSZ+eOaBdntopP8Ncks4QX3ZjslYlDHcBlIwfjSpmMQDlshQL+o+4kY9qwSIjR
jxPdG3Oc3ydC1zdXKiuBMpnABbyPBzGR6p8ayZeFLhigPQsYiWjku6To4ZdFQjejTgk1DldNaNlp
R3ixYuuef4XUdjArGQVTWyYRqTI7u1zrVUZXtI31Zcl4aFINjHNNAQ+WCADWcVrockcOiTtPUhN6
pJgSPm6q8NMQY/Qsb/s8sP6vrG440vZuo18CPVAbQJg6WMYy9u+gW0Eye1pvppZo02HCjjLgKZKE
NTucdmZye1sBWdAiudqBKmIXGy+rAudEbAp61m7fyBg346JWZdhyJyxF+1hB0II8g3oqlt37thLx
83Cg4szUUJ/JmjIJRVg6tNsWe2YVFbce2D34IFTS1aZdxqCG5YiKnUXKQzohb1LiWxEYnkExiM7s
vzkXRHsqTOSvc+DR+xrYr2G13OlcsbgSUgodgO/NCgV5aUpOWKMk1NC6CI9Z9UFn9zIlRsvL20Cr
xQs8ObpGsj8vJ/8tEjBuV3B0LnDtPBeSymdv95vlYHjhb7gpcyVheFSLjDZCdS58eQNErkAxgQAc
bwZyGgZx7IGrtlpx6h4HeFyfuf1ybFsxLYcZdSuoiJmdekkB5U10gLyptIJ5ohnTMird3j63A8Ul
NIauawPvaHhnibXxHihbQqLTd6Ka57lJNM+3FIXImpb8T8bTCZk/b3z+L+cQDTt7ZiVbZgKv+kq0
6SK8LTe2/r5lyz92M9arShmPzozuR4xl88Gju4hoi71optu7R41YB9v1rEPduQq02x2KbB7Rhpsh
/yMIuu8IldqLP6azJ70SPxBVe3goysWJK5Q6srpUrNApNWIJJyRxCDSXY+iXZNrJXE0dI8C8DS2y
p2ebgOL2A3tVi6PkLH+rD2NG96XIwe7Jt5RYldytLFhpadZJ4cq7TxioijSJ3E38Yw6JS7IqS0qS
jyoZD7yxvUsoQH1u6Ls7jn0EADMLeBpPydB2yoHbirQrw7nHtKL6sR3cNJZd1XzgA8CMpe8c2+cW
YwXj4HRCpm9hSdPJqnzhl1TU6EdlgEzDj+c85scC1OfGpMZqUsj9O71HmDCTSeNvV6P79gcJRmrb
eqE8Yv6izmkQn4AwvH0NJpJRlme4rDdkS7hBR4928xvK75j4k+bC+aMTWJW21nyUBaUilYaux6SC
4X/3SBvTMAXzssUhmlEoiCUTcnIjjU10llwU4vp+PFHJjNjqo28M+NBApB8dkvRbw+wxZo0nBk2H
49yLm/+IPLDMJ5+6JUEbTsOoIFavD5oZ6c27D4Pas7aAGL3bixjlng9q4eXxwGn5Bt+6tL3ZkkNd
vw0VbtzD7wA5YF5yrBLgcA6NToZRbFLQrlCeR+cQBlLx6f328i9NJPJX/3rn3nX8HDeXfxQdoJs2
nLqFrHoBpZ4PqqLJxWltY7ce3qFmEZVxTrtAwYCsPFc+2tItXna7VWXUSCm9tQCmkPavgfEqKO2Q
KpQsfV9qk9CnxHM0YceaCM2OSIeRte+hHhOtCV0QY/umXHqp4YvIbkk3Tp+c10+Y2qDYSD6GAERx
WaKuzrr4e2kIp4uXMzQaNWt2mOsfDjAamPu0SR3CKd0Rbbp+hKE7jELNyxXiMFf9u8F6i4Fl1Bca
fjNE2QrOPf79spzIZINPGEU2tSOfG+S0Mztw7a1T6Wk3tTkWxepykJrjbX5IvO41Bvj73sYJ1Lmc
aLTfnpuDZmuKjaM7DR1l1dEHALYdC8ixJzcVzZEjiexhDUpwzSSIgVRzmb9O1ua/V+MruyIsbuOu
f4KqWwdxhYLfHyJftzt6MEZNtcetb8OqKWxJobVFc1RmW+BkQ8hFyNIe2nB6cL8ic2FEvWv0c4mU
mDifQjDn2HnBoPIRI/0G3Up2w4Qfd98Hzpxv3lQE/fHr98lbWuThX4zmVpUl9JTjNBmMpuuQdxlR
1nDE0+V2GoNzpMBXtnrJVmAEN/1pVDRkykFEAUOp5/brzN4Ev8lxRQ0g45sNliR4NccqKAXkAoHk
wf6kpZNyJem+Ynf/3uV19H3uxEYVvdcWp7SyQgHYaQ/cD59HJLT+I40fxB+thkD6tlnD+woANj19
eD4NDt8C86Tm6LhJ0LOIhLDJ152vsEjVSbGu8g5OUt1OlY4oVbb+yjjUcgrKK/XdGjW4jAadg91q
x2L145EJ5IMNk9qZX78JYyutkxV/aACQbfzA6ae5H3wRkq+pabVxZxunYHe2etBQNPfd9v5tv6c5
cyTiutUIG5BRj3rfm7BQRLBZr0Qqhpa3Wp4V/JDCAQ3V0xg4SfGhsLQPZznj0FkuGO+2nE/QdKgt
35Kxh8WsvtcwR+jIeQ3PH/2Byypjp+zBiCZB1Q7dmeOVQ/IPt6YimZpLABddFEg4qpCODqH+s1+X
dKJKA8rJSHJ5ZhZr6SlspwEosUeA5bX351qTga5jjE+2yRc6bTja+pCZlgHA+GWgp7Gt8LxNEBS5
7Xg5pszulNkEwiXSrjhtAabAaNTakGoPXy1yTgNJhhAaVsvdtwmJeNPiUErYXRFE+5nBC9qNBvRP
tlNSAy7NZ8eTpzOPRY5DYHu99SfigD7zycDL9NDbhCWpRxMQK5DV33SMz75McBQItotN7a2TUyAA
Lj2aBf0LKmiIj604VUofLXfeP7QBVCMD73n+/RWVz5o+S0/tEPXbte8iamlR7IJ81TaFOK/1rIGh
AKALj7wk+fRU3DgigMsDYj71bDEf/+z7W9Dur+2kfiJXsenGAwymo8FiJPvWapMjtNNwUYDOsXv5
XW/6RF8q2sgsctfM4OxEPXxboDpZ3/uf8d9rbA61xtJQhMFCBFaRIUHow6NWBFMQGR2MvE3mVlGN
OUo0QklmW7g1xgfUKQec0kwXpF3xxcH/NkZoMWiC/eF8k+8a+EkmVHAfsOwYa/D5B5n0q2sm2SJV
VQ0h84Iviro2D10p/I4RanMdTqLNzgCMwlSL9+hFoYIv8loj0xoiy/8CuwVslRexeqWa49xxaVdF
MHMDXCM6uJE9FQ1PtwcQbwIrGs85X3nnIYedvKCYew1zkINRMMRvI4B+1TgIzp12EVXzCzLSnoHc
XONqsf7rl1kX9JtydUqh7bTNyI2L8FDATQm+ZjELNpOwC2nP+lsxiHwYkY5Nffx4AoF6U4vPjCoQ
sPKC960jaixX+7Uh0PmvlywbUXB0D7G92UXpQd4upZNpe4inIzUm6aRPk1khVc1OZUzNQWBbkmHH
fVNe8Ae+//b2R9BAXF2RpXTn8ryKALJc0++72e4TsTw5hT1TcQR7Kehg6dkksk5emPfEhCsOOmKM
IpAErD2CGR4SUYse7ZEttfaiqoZGAMbkzCdf8CnJgnraYFGJ6ZpF8mJoki5s8oeREG/+IieG3XIr
YxSiNJNWttEYwT4eaZt3ZKON2ik5O5xrXr9b5LQZwExg81NNdgsIUkf/qxOUY41LFEM6kbXmlIdz
tiFa/W3/tNtZmIKNPM0fU/0hCaOzYbUaStPaCrFm5yQIojkv/PcLk5PdmvPxXQyw8UL2K5bUbXZk
rQ9ck7zuJmPmoUc4+UfYSqi/V4i+qJGMtkyeyfnWHEAjb1WcOWzidML0qDNsgQ72qehueW13o8ws
WvzLDfdfuUADB9nQo63mAqApcuWlE4YqC6SyYEis790+WMl/Q7Yj+bZ1ANQp0ywUe8L1nXYmdLXg
BBG8Xp4j6DtLxryNkcUFWdnKNqPipI6TAH5LHswl86XZeAS5AijCRre6DHaKLeZe/34mODkcNXlw
jP99TSjcwNMI9XqtyaUlQZ9T+Otxdat/KyIv91eCcCEw7Z5O1p7ErvcphKA1mEDQcOJVvHiSYFdU
WenWwwxgBAW2tTh8r43WM7fFfT8D4/VaCsphg/sjILFmFcECfVuaxiyK7tMkIS092iS8p0612toU
OM+bjcdJA+1QvJL5FrhlLnbM7bzvq1tN9PPIPPfrfB+q4GAeGo6Qv0pd+kJgysMeT6l/J44clDsV
NJjjJ36XljXjJUBfq7OU+EJu0eZR5i8Uu6rD28De40bFjwSE+LJO5M35kOVI/vP4DZsmVmsMXbvK
tHX2amRnZhCkVEKPOu6Qo5OewaDTgCsn/4V8aTz36jF9qWr54RIhWDKVAk1QadyBm7BY/Q89F5Lj
UOd6qXgFACZRK0wgdi1oamWNCi4Z2zw9w2799GmW4f23VsEmwCdClZheskXM9ZDgALoGv7ICuWqi
q/GhJFVk3Pa3Y+CL1+Vrx2KNsDk0KSIl7gEpzu0E4DIn47qPyHr6oiYK8MAkh5CrGbSw3lNs8Xl4
fn0ZS8JYl9R4dmHH7U/ruH1waDaLVHK+oCY/Gli+Sscw583LC8oklO2bpg24gntvYJtOsPQIGNV9
Nl6QBZr5iTP+KBF22ZpYhlgdTaZbMLKHZ+HuJqqlJsNRNd9ShPXUCNeSkOiepvxzpFJKb9TnnYtf
0lcD9IvilzDUVD+CWBfgyRTCCFpLUC3FIsKT2PL28MhGPaTPSXIreTE+0K5Hct09SM62k0z4x4p7
J4HH5PVDNs2WHOIpt3O6XdixQPcEH+It7QdadbLXwpjDf/mZG04TNuRXdB+kHQaBz+UOKuQppNWM
ahizqs3TGDVWgbSrxn5hHoBVyB6Ec1RIeFZOO3QDHNNcFQKP/HGsZbD/wigfPzL4pYJ7fwcGQv9s
VVd57cs84kCX7lnSJVc6Gu0Xy8Xcg+T8j3Ak9/2W6Ga6Y2HoWv+SmkibnS2yidXSitYyAJwx3zTZ
S65FwebL78yKKCV3CJtJpgrrjFFTVTc9sQYjpalctePAexarjPtt3q+13EAm5OZETU8Ju18fVIAi
fv1/38cWH9llp+r2jUKaVjG84y5JtIwYWOmHWlugm693LB3v80yuAyT7WwSMOBtmQm3R1JFOd4O9
p2S8o6OSQbJrPNcnSopNUlovWKr4tQNn5vBAFnypDcm5G2vLTvuMIuSYM3MI0Q5728V3UIVQKlTl
vLtuw/v1zJiYNJ5j2O6zL6SsGRb+gtPgzOf6FBE+Q1YNZR62jrnYL5QS5ac6WV4EnErkImzJyvRa
QYHTQcHuhCMZsvhlRJj2zd/tOzGU1dZk8obpXeWc4xVKZvpxQ3lpNgRbSENGAy/UtRrDzuO0bPjG
I4ChPpDOUM5WeiGZMewklTyqhTTwaMuJoxZetQcqqDy7inLLc0zmM7ja5wziJSqXMoQuR31D76Ti
kpMZH6aM1Zfd+VEznst4kcuNIpwquIYzzD2mpnhRllE1QTaXrpdvp2fDyfKXp0xALwzkFsXXAW1Q
gmEszBCVKcOlVBt9G1Fdj4mbqjpoqDwqhC5qnFMx5todk6B0ztTGFn9mnk7JriLfvAQc/5DOCOj5
PStkvMw/fF5S0cPPr2v/GtoBMx9+my7WVF9PO8B2eDKrsqBghBDrbiILa+DsxymJ5US7oiVWGrBp
kQh/VdXBLaxF6z1gYy+QKRwEw7i6/kuiPjJ+k/Av7VYrRA1aHarfwd3LDGXtBIw2KfcviUclgbIz
Q6/uyt1ucyFhiwSVCtHGvVaTBaFNVTiAPl/5y0yG/kX27aLl3ke1t85Snlzio0VRT6IsgfsE4mBs
q5UPa6cAoE3JZa/AisEqnYwOnJ71OQTY2GkEQOJCuW9wrUV0apP+XqMTUgC2x9oPlj9Xamsd+hTU
pJmpSFnGG4J606WdsTaaN0DwsyNuRGY6qb9wUpkx4JSQtGDAxWyG2ZUm0WkzJ83DHTI83Gub6ziX
EwA4JIQr05EePe53MrxTPuFJSNjXnAwPcFjJ3TWVGteRz7jKp/RkTxMgfw6k9TwSV34hHO0RkWg0
0bnXzyqvzV6ozU0iNJOOV3lCaL/EQ6oTLV8EhWfcyYPTaW7lDd8Yy8QPrQL1losiddUOuVA+onks
RVk9FdvlTeQglEV8MFUIN1CItKvQ0bTPEFwY5wve2rSOwbqha5S5ocDA0niDepJ2yjrSZO6qJlKz
1xq4PquPxoeFgqeKM6a8tVeiPZRoiklImCl1JpzByvA7MzrzJH7ZtLQKDdkUA4ZkSzYKRXaQ0Xn6
0S1mcM94RzgMNLyis54ZuMBNLX7XYoZ3XrwWJgtzjMyJYnGIqXFfvD8YA6x7+fFGCtWeQLxFBoJs
Y/aBaUtlEPpbtMnj+OfjtYTcQRhiK+keKK13jdIpiPSYXXvYSwAfQ2juCVWjcUuVl2Fr70S05sy0
7TCojFwLR+9WTIu/1E+BjbtmQAD2wFhRUfl/Z8fmIx6QW38f82Ar7FmZAdXZzrX+7rZg1/Cn2yCK
RKGRBdWLDeZXGUfIas4pA1/rQJh5OPOQLnP6IdUmC3T1RAqem0iREilEnFoBJY/81a+SJ4/fPIT5
HXyg/+kXKJun9N5j3BOm9y0Fws563cRMQfIDPct152qQpxj+wgEl02ZZM+kRWw62arx0RmyHkITN
rFK9K4gWhEGi566qKIEXDHf1EewFTXWxmsprI1qmG6aF1Qnw77jCcId7+TPLOt8nNcAMWVJ7MYg+
oc1UalxA/HfKu9hsGzPJ6+FP8DP7Om9ZBr1GxazB0W5AnJv2r3IyUdklveXGWAWdDGfCgf5/z5VG
YHWCdtgYCRmel2s5Pwi9g8YOi6wjX7Tyz4C4VDQilgK4DgMMqCAo5c6TRCd71sRh2j4vFhIMEKq8
Spi/GyaVvPToI6Qvm7AKl+20yauSvi7yRnL4RbrfZwnixtUN2Rzbv3jOCeQ0332JqLvEvr9VRl3W
G1mGIv8EkjEzC2DYeWAfXL/Smyp/ihyh1lssboZ7nqR9hsCGrQpZq//SNRdsgCAXR/R8qomBLfha
kQr8iP0mFVqzEKzwbSe/EcwidPffscg6If2REzQd2qik/R7NehXqCYd2GcLsFUVIrS+Bil59aKbw
eXoVL8xo+i0M9KjffmM/sSZGLWSQalTj9Ft62wAUjBtD1yGN/3TjZOoCMTsmXexTT7a0Mg1ck/if
R2PcDqS1+2VDYjq9V9GxJ6n05Ldarg3qdD64ahY6wCuKUh7Nh57a2VnlMNBFTrQSvD5Vz5Llz6pT
YS82485sGpp1ifSC2eE/x5SCjOPmJx8VceGQ6lqKQ8/HjfXUVQq3B0HPozqr3kUc5djXyOlVtYax
982SPNM4UE7qSpxSZMOwMNVYVbqzcUKoKeQ9i4gEB60a0gJod7FwLGquv8CCtt92XJ+ErQ0B0HdO
WzuF4Dt5HJFxXkGVrzu6YXHukXHRba7YU+likgVHdn/PLY2Nnuzz56DkEUlyKx8XP9gjEoHUUdax
doub9IEjXm3K6+SVqdjGr3Cc84QP9KP44s8m22UaV3KfVLWprRCBxIF157MD6M+6hL/ANMknRB2e
jhVvRkwcap6LXXFs7kNaxeDW3LltNrrnZHxtSGeey3ttA+EH14D4+PFbkfEnv0/F4ivL5rI8Yrkp
ApFXyA9VY6kVvjRwktphodqsD6WEpJcZ9boczWxcWgARQtTeljwqYrcx6jyyQDv1QYU5mbZEB047
gmsEa8b0m7bW4ZhlLEVvwTWagYbDunRyfl5Mrio1bGg7iWjUQfDiK00YJOro3FlLCEza/FCMFnbE
ihicQf0IIUR21GkhikUG/F8R+RCW+1WgsEWNsE8BryrZqFHaEtJuiSUmmzqKAbrxOunN9GJwLTUP
0f6oVEP8MunOiAc7rukbzwMttOJItQtGJmjQoFqMHKrk+MZGqKmEGMZQzSKUNRlmrX/oItWWYKKL
FIluf7i39n41U8Be0Fck6msTttq4l5KdiG9QLarsLBqA14jLXBOf2pGrdaGpfqvX0QM+zeleLzOF
iuAJNmkBHfPKgbnyO7lwXXne4oP5HODOuV1yu/onRlNyIS/URMpZqK5hIhAL8W29YyVci+zaKEvV
D5tuBE/yovjfO7GZj/jHaOlr7/BiYGeCqzbWAlQh9gksYouxMQEm4LDtz8cLuFpDSW7jv6h8qmEP
IzMGhflUsSHnjuk7ZwZVDKCctqS4BryGueR5ksZb3EiqvlsLvDTRM6MhI/Q94C/vX06IXAlkNX7k
xKIMcdipd00MFqQcoql5dBbxk9FOWebZtlMdllAE2/vHWlPEdFOEbb6ntCDOUPyyrwdn4Yp3Y7Ja
s4m8/SXhfu9OM2WgqsdVxZ4JbKgQJpKDTF57CQQw80reBNRWiAlO+rKtlWdSjydMZ88T2J3JRZrd
1z1khEhUJTt9fjsW5wgFd81HyM4yO7Lo80FxYl+3ZW72EM93MSdDHV0LBexg0XiULKdGSF+OIotk
yyCMw5VgAQ/hJlA2bI6t3I0cCUcJlCtCBL9Xg44XDoQ9XgveAWzdq0ppdBwSOnfm+G0IY+ObB8dz
St7YTRBnLYDFh0F23UAYYMlkkIV9KbRcweiZBLu2MtZGLDA4j7grHuI8k+mymsyVWo7CijRo2Pk0
IAgEjRGHSEGNYnJ5j6xzQc2/ofKYC0h4elA1md+reiMvg8GiwIxPS1+boNAjXhrOJlYdCx5UuOqx
CsrE05LU5UKWTBFFaSfl4xCHs+/Pb/+IrcFfWqlS36cXMDeJp6b8XWH794c+Q3bR6gY4hRwiZzXT
McFjhjVxkLbniah0O0htb17TwxrCzdcDesgiPdlN5gbfCroikbxYXG92INldJX7iarXpBTi9BnbT
LNV76qlEsSwlMI7ERJGViSUByeJ54GdZhKi7XuzA5JE4bOP3w4/0UzYbekk6ha9Cb8+KXJHagn7z
8Pe1DXVGNKLvIlcNimF//g7Uwc0AD/9rx3ED7BsNJQGQ06oMfedyiETErK5MpYemOyE980RX4aR8
Qe96iD0MH6mfM1xh7+lPGAtipxLBJROYHIF+iBz6lBo5bpBEaYSsEWkgJ04DO+6iiwTLeNfxYZTi
IHn8ThIruSYOsQsODmcC7GBUr2ELLbVNMah862dJqNUE8vocM6YENQ+7o+Qt6mimurtwJIpVZAae
Li5ls9jjaZNCabcbSWTn8kj7rCFVTXu8+48MsjTTDyTEC03eJ043WrPYTcmqjCC3IXW5QodK7Psh
u9xEDwPDh1LSHO22fYKpb3sK+b7OzXhRdJbR0l8JeZlgv06ccJzd5QkCu9MwsqZxY01TYT5XCwdV
hBWZ+/QmDC4vi81KPMgBkx6RoXp6E7+WHA82pyaiTBZXyJq/B4wcXEFaJhIKUXkN8aXAIFGbcW4t
+dzmFR/liLgttuHUwkngJU7xw6boI9eJuYvjZnihaShYco4Zn32mh5s4drUUkwGM1ZGvdylfcZPK
FT6BQhGHE0V1oHny2HiiQP1AfvzDvAtMTVpqsNehlyvIxnrR0lhub967Z3H/XGqqeskUiyuXBtp0
nd1Tci1SQpaMV5qwiXPo5+z0OO6f7xdIMXym0dw0tgppmoOn1f/7WXDfYF9x0Oc+05+GbPzGwJHU
+4zuGCY/TPa2XKiWkjSSOCuRqyKJ/6kIQvT4yuPOfpohmK8nmx65Rkzf1JXZbkiDHQ2GK+A57y2Q
5CM0NSoCYQu6O1Yw0t3XANPrwlH13azYdHNN3kdic9g8/h8ik5qxfv/5SmI4VewwP1lBy44RTcGN
dKdILs0XuebNDZCIHLaA8SJaJPNKYTu6CjhlwuQIIl3WOtMfRa4IRLYf5EUXHIz/QbykDlI3a2rJ
4819fQGCi0pSh3QXI/mtI55acqQK4HnIJJ9RhCMZk4bWLy85O6NtNwhipJug4ayWEIIFXUOE3D+q
5eBAS75fPhgE3YqKzO76KnFYLD29sFDIcdlZKCUYFIYn7ZnvoqnyvOK/TJpPCR9j4RVJ/W0OJrgY
7jxTW63+Dl2nrmB953dbeRNKj4K/2rI8Zpq+Q4vLl/NlGw6GF11UgMJOvi6/6tSe+cPWG7Z/0GJe
HQRQCYfP7fL3sLoVeo1Zo7tUOoRn2hBOdWpCCznstMN//QyFuhwBcm6NRb33IxcWh82WrNg605oj
3LPAazz2jxypUz4L4zxG5WSviEnf7HmJi1zJShnv7nevI1KjfCHbZ9bZzKY2fVr6tmZoO8M7iK7b
oK+jiNkNuNRDxzmURoEfpOsGBrvUMWnjit8eZLPW93g70rQ79Jb+SfAj1w3P94EZ68pLl9NVGril
yscofNeNX/26xWhVi6h0ejjfgLx6dT7XrZN79EWxcMTX+fivAc8CCYWIKL3YAMSY8XkCBWSIPdkR
NVwoFJ8kWt8LQ6RJNxCXqXSqNcBKPARXHGdhRAEK2ykfYxlwc30+csmGWO4xhW2UeVQ0VErm1VDE
PDmosZ/t72CRSOhq82FUEcfsJekFYtp9+7ScFas+MlB33Y+DTj2ocRfx7GmovxeuC8hqvPDkQROb
3pdAxzuqv4FGrd5S6xMobq220rhWzIipr7o5EjAx1t1wfrmY6ImgPRWymzgbFoGGXOBpm1+p8nCd
cdW9F0zPLzE7JhG8gh19oLuSQQhU+hlma51fTJ91MUfCFPwx0AEW9UyOS+iRXRpwmR3NIYOpZ1Fy
kMDc+OVM0P/ZPnaidftPsLVJ5IB9kYUoL/z1mN5V30WnUXgNU2cVrHzEYAB7VT2clX2RInuYh69Z
4ROt3eXlTnAPl1aMKyf/A6slURrDNzgRuHRZLqvNTQefNVJTfFavsdKQEOSb6FY80HBrRx+uWYCH
Z9LhkBf1gz9Bnqm7E+notDzERlqRwBSmd/XVUNjHsgdKy86dMt+/clCL+Sc7c9Ih8xu90aMtsC+r
V1QnIDJpqrRtHk8+nJwVseFoXq8qQUCVTaR4SZgDPyhUhLu9Y4lSv6KNaKnpV4OeyFIkHadJi0xU
bVDFIQHrn+//0RwNlXZu/US2z7G/uURfu5RzULBFr0yR532jaHD7FDZwsOa4Ci6vT1rEt4+piRnA
Y+OgLXRz3tmWv0++O3gYiDu7zQm9djRpQQQBBVj83ckCkRbLbMEDzzuFhBi7X46tnV0GTyD57tk8
6tBiQaWbZoByWUCe7MVpsYJREFHMlwaAPTtRTKByRkb519ZKYkfujh9sgl98VIBgh+oYDs9D1x46
1SxiqvZTs6fxoFZbrZSgeIfLVqkJl/KSQ5nVw8KXfn+ERXqEYTUkhvUfn/Xv0bmDW9BPOjnEP2jE
+7Er+PAPVTHGLBV9JiVCtzEUtXair/KNY+HxaOD0a/M5HpFkrSYMXmMtSz9rt9qIRIXGZoFsHSIi
R5deA/2GGzWCepk432MLgW/1pz0YcDt1SE7yiB6a1emr4zlgt/1OTjGJ2uc7UhV51Rc0ZONtCm4p
nfuE5c5B2QFiXF4r15ynfo7BxZUqLEN/xxtFgAkfmiRJ8pbngFu7HWtH4LB5EMgR2T3iWfJBaA9u
iJ/ScLNPS00qpNsIHrEs2duTfxyLXsbq3u1E5SRItzlFE6MK/VvP1y/Kjn7Vz4iASZrokxS+8tCj
W2HaADemL+qFb2saax9wA6ybXiNHkb0q3jUO5+19ZFVQpvvYLfo8RXu5iaSjKCZMZtD5xSVDuc/F
o1Pomd3ju4rdJgVeeyitGC6SU3o9v7kjOMEg5h8CebRzLZHnH0RwOaDMrQ4JOcAjmYvIZl4NAYww
cea/vhb9qPD74V17zsS/gOYvGaSpwz7jzVLBsmQofB3GyxccEXso4PEUJEnkENmtMSS4YXcEHMJl
qaKXYFzTeZonNB5tPawzFr1szSfSNEnZENTxWEJsvFZPyz77GnXq4ffU7eR3DFY7puKapcX7ThX6
JxY7+vLP0Decbm2M4c6ElA0BfQiHcHS6wqWhHfqOcBwClRZywz1rile0cEKJKn77s6sqs2MAgcu9
VhLRXvzvSzAPIovB7BKb2LXjGOsRqGMzDFmhKZU3uCP90MEjCHkQpVj5QSOBGZf+ssOGyib+DN4D
jcKdDd12KgArabj62Tnz0My6IjMYtwnNonAUNya67NZ1AUQvJ86jJOL52/BbqlA9C8R+1sPFKPRC
5K2Ch6jeafeSoXUSr21rCHCLK8qXuDCQCzM0rYOOTLoq1yULyB2tOG7Ha2mboH7uU+uJFCdDpeHb
Qu3hdK1DDQqpLcKdgiBc6aBYU/vA4HzoQogMsx35HZ4jL8xrsd1f4gUAeRkkMtPgUpDAaMwmKRHb
1Cnb0yneWvdUr58dmJMp8CJcc8uKm53kM3jLV8BVujeOTq99p5NdULF6iljqxwcLs5fNuMNBA3bd
xP1qjMzjpt1UNOKzJazHiCWvR6CM2NcbxDgLkLT1IEsaB1KTck9FLQhrKbFuc2g9cXYmcD5DK7MK
yvTlXZaO0eXzR0sZ46Cio0WGmHGHBbRGUV/2uaw07dzXfqdF4DCh9c4fXWG8eF9ApTPZLxQvG4IH
SYKiOJXAHfBjt9P7OGOHU4bH5cI3C5yu5zK8OGtsgZnCfrytwOOFwqbWAqcP+2DsMa03zM/a+3dC
9EUdfi6ZCC1z9ZvtfIZ7GCKLL3nnjZLM5HmnsbDsKLhM8K+un3VjUYie9vaHWZxCHKRKbbCZKtY8
wiJD/9PTyc3xcVqCKkh556Hy4xoRA/Anqs9HVHcsn/SIx0DaLBIlOxTzq8X+7RNZHs/eNVxodGfM
VEpXnuqwuOLjyCRK1mTy2h4o967I466/Q9Nit65taQ+/nqkOvsQzvaBv+n4JNWUyoJmaT7Ji3GyF
XOQ25q+5kTaZ4wlaEoETflqB6N4coo+2dk3L9cHj+wSW/3+hL4btfIQXzGYlv8S6blfrW9YzEE1p
IxHTRYvzyROeoP0mDVYpflsaRdx5VDv/aJqgfedjrri6UXIAbuEtoXLVPaTsxlo8uUqhPk2xgyjF
Cnex5cWiKjEPjpM0Rn8xO2f6nF849GlcZDydEuA1Kx0WEI1haOvxhMItKL1VNBQR97tnRlVd3Vyy
pdNEbBo4fg0qA4mDjqNIT7FwmcvHLLuYfNZXOKRYpKFW/QHDzUiusH+lJipCtSzTl7W1ZL6dZ8Dm
WZwvD894BbXRmZgGd77koebziuweJTpeSooYoVpX8Kmk6Qk+Jn06x/HhuHlL0IFYu8NdwBfnl6U6
Vg/jLHuAo/kcqH1UuwY4E+ZSrYFTtDEms1+agBwzGOYKo+50wKduGYc2DaKlBSLBS3ivgvRnoZmu
cfoXZZxoo/CkeW69wNfBdB18ZJFqlXHaGnOJ2ElCIFwyo8nf+EVxmQFV71rNzoHb7zeINe92l6s2
RpHlWbiw5emMZKl7QkW9HwQ5CPMDiVh/xslfCYvLB7Cr8FFgmWcZl/tBCn0pAMEhgqbmarukXCag
aPDZ0CoEAsBvHRThQ/JCNk6O/4gqDWW8W/kVXBIEzouC+IGOjurEIwRAKm+TLy/6ArSHicMCxLoH
pwEQ3yEj35WYMqD8a7yzmIl2mEXfFRkAtDBB9QrowBe0aNZshxGE35Uej3Ce4jsttJzDDhQwoKuX
sRSRvv/7arH+eBseB9ZiMZtH9UegRKufh8Jo+kNvzl7eZkYCpTAy0xtB7GIJEeKOEjS2peH43+0q
ptnG/Q5JrFVuCimbSNzam5U8O6S8LeJbhDxt6wZARW8mCJlA5z+nxToaTgSFe24ZJlA+NMiVx0tA
LwU1R/SyO1DIbaCO3bkl7H2vzVvPmkly8P2eOgJwneJhohSK8O0Y4CiYL9JMIl3MaGqWAZHUyvZ5
jK8TbfoDLCl2C9omRFAerPQs5YsRWZy/XTYweI6eEQkuiyzSz2QHUcK5P69p4uzH55DwwAS8O6Uz
aHIcq7hz8RgsNEMr5sHwl6P9UH/trj5IcHxavs9RNZ2BHCzJJ+00gNNGhuLltegndAkxoFZ6rrA0
6XiLQKURxu/43EQnB89b4Mpmp03zQpfldSIt5hvQ0ZaGUvgKb5GxIlCnEZlJnZJEtktbYhsBPEIv
61zucxqR6v3moFDo+3pc7AMO8rbOOr+ZRUakE8butO/hqmu7ytVsQAAX8Kj9SeovYxCjYZ3uJHZk
AD4Wh4M6hJa1cjU1ZNxt+qOp5i/u05U7xh7Ly/SmluNGrCKLoWOG1qwcSaPj2MmPuiJUrEUeQLIX
I8rR/VLgI7Z73QteYOC6B/UVeLg/LKOUI+ChewG1fMi2N2z7mH2TVb4X7tzq+Ugbc0k3Lgp7KyNz
5l634llQrnivuC2M1fJNhMBNh7ydAHMnUEqaed93GVjEnyPBMtIBDI5sfmPGeLdHYTzuzzOaXjCa
C9Zyp72fjaVf4Lm9PXROuQGT185I/9aB5bRYnkCN852PYrfJT9+afnwVTVg/IswD17SH8ubk9KlG
Uanl5MtJqgkMmdZnJ/WKLmbQ960zhFOH/IkHdz1v7AjwTTglIUYjc89Fze80rlBxi0g45gbYOFas
a0cn2jXQEivshFt39GrtF32upl9+xfXI09uCbjxfl2efdww4uWEbBb1vCzQPbD7FIfxRGLs2E181
nu5kVQrPOSpgUtRr2QBKOVzE3/uqtf7IQ0XPYmoNBR0OdG3p/eUZnDQPRjf2rZxVaeygVmciIwRd
Al0HVQ2VI8L+S+n04k70eTp+W0N7O+D+wNBklrmkgnhrNeyyvXJdkjIPrdz/26S/CJHI/fokKdAT
GSURxP2QutjLnf9F2YJyS/zSW6UeG7J0+6z7lFD0xrIs24EkIrHb5BSArLdUl7/91NTwUElUx2V3
OFRFshAfFNBdnJh4uMEX6lAzuFI4gInL/qh3iD5kx15V6wEleZ8ZR00o4MY4gkoyytGPfCG+392P
Kgo8GtLi7Bc4ik9pfzOBX4un6HALizfkLlDfgsz6IW5rO7pvafkXE4pAlcxod9BdDwj4WLIbLRvE
p9GaSc6FQiidnJ3F8X1R+olh2NLCylXxrXRwkbhsUDw8/JD3xVZwG7BHc4zxujQYFQEX8lbLHFCk
ddgcYuBNErMpbuSNVydfI9hr5yEc70F70WoZLyXbTvptEivvmDbHCL6UGAfCornaP1YFr1oPC5+k
UZqaV/Wsy5BRnhlxa9r3bHtfWtVU2+WSG4QIdBzv+S5Ad4pDNeBaaQ3vAZ+EDsh1BYgGzL13HmfD
ilPnvBarPM+2B0HUAySKwG3CJusTZ6hURnp55y0UpC7KKKKUK0j07Iyfe/T1oYLVLOaLQLsjEnL9
lkMj/shTXz1gvZ7wZJ/LyVyoKoDtHRZnDkvfUXv+NPgiBrUXS634tUr16FX8kg2JkrGLuzrd5XAt
aSUrModWrU6KBeoR1PpMmckZzc9awWUvwZuJtG3ZywZYa4iQZzhuawB/Dd8rwHf9TYkeyQBDDPkD
E3Opdgq43Y5LfpidQSvhEoJ9CLiv8x3QZ3gTBBg9vkIzCAkn0MNziyOQMEdvP0NIL75lcEH9Jb7X
YW/eHLBC74S7ToR+sIH5g5+VrfNoVNAcSy723vLVMgqH7SjXpi8EO668Tl8cRP3IVNRgyGJ63EJW
HQm7J54ZV3RamUwT9v5JNRpp/p04DyDVhNy+WzsIE0kRWd5ppHC9JvoJwnUsC4Hf40oxyeD72Rl7
zXC9S/R1s6+VrczJAGM3pXdryZNNlvgABw+FiM/QeBmAWnPyHKWdzFzoxcBgGcnEDXbjoLi7myML
vPNum8Mo3AW57Zix24jnChDh+dOyYbNx1MY4z7ukQj2zc/Cp/A6LbvKLb1TxNuQrckkrXYvSzn19
1RXagZ+g/DgSFEWRaNbM/YWgxJ4NcDi3q3WN2PEEYd50tYqhA8Er4Lv+DAd5Gc1P5mpQJklFdB0Z
xrT5coQUj/+ON4aFrIcz/Q/SMxc6eHmAnto1mOm9ck/X3CPYmXvRfIJE7tje+t0GIecfUXKuSNaR
6HwqLovHPKJFcabHgYNRHSL6D++vspxWeLIjFmIj0J6VSLf5hfXXrf03/y2TqNcU45yje1NmEVBW
5nGa0lFE5gds0F7tww7HX/o0JI1j2EAzBLR5DGaQ7++ORFUrqqRYzA4Z6DpkN0oc+qFU2HrRJKBb
rR6aMTzjZO8/bybWhGSkWEIdEkwXx88yo38EiKDCeGDGhFEAdC4RvYAP+GthISDp0ggcUm17O+LC
vhStBz4d9s8cJoxNXJbqxGeXxa9cgEQ9XfTBY3V5sJfDqn/LbBX7ZQUoU26xDXIJdLkVse8m7/lG
OLgHIpmKm3L8grR0LaT5rJ7HKJfyy/714uj2Boe9VJbvnEbI7hONOx3XCqQELJkiKsITLZgWnwTt
KpCl4yAYwHDvpoH2UToSHeg8Hy0LkK4hPT3ZRf3ygSikSN4AxEC7KcsZUxmhdmC9vRcPn5ccwea3
yvula8MY/SM06B4aV4EIcE7ssBBzbdxY2y5mieTGNZfWfW7mly30Hx2EcdRHwFoHo8Ek81g4VCZb
F3b2W+k2RdCNNStxN1JqnDOSDEmJ9tmim/KQhSacSxXTF7Pd9kFlnpgz0sZJBZPjZ8xgQh6KIVQ8
b6gD9gclsQF7ad6BFsGuHcPuHmVqkZdkwsYjzM/3ZIMMQRscCIjANuxg6f8vb3IqJ5JkYnUdG5ME
lpe1gLS5L9diS2j7NaUmyzElXSSXhYqwBK8jy9k+TlvTQRmzu+82AxZ58PWi8gIWwN8b+g+qU9Ji
CdOTOOx4VkeRyhzuGTFsnrV293k3bCvym3Fyz29QqwKZ9Z9PPocZi4/PHbqCgCysehiGFo2lsH4Q
R4/EK6OOwj1r45vDuKzG36bTJgcGl+YUeof8hjnHLRw2WhSM50hahRjUN24H0GX2HCQU8lQX5YTU
bGFDnCYtE3RACSFxnOnrBKKZ5sbfawdlX0VvVA5QwSDfx+zjM7noji7BTIbGRdpYsCtw7/QaWAel
AltWjYM4XiYAXwV8FHpjKVAr0TgBRYtKbhAYcIUR/fDZAQD8Y6LuU0Uyz7fp8gmF5E2RQn5l5jvb
l8Ec4GJ9rXrWEdxg8gqa6avPKa9l3fgXUyY+CWQMo4O9srFWJVIJlnPncYFNhvsxjlky613iwYYe
hJMvmkK+OLEkkzWoZu0M17uCgRZneXjS/RAf0tmp0aKpDMF8tM2lYhXux+UAlWuXO92pAWMmXvZY
QAyvAKdnfu1SGUM1SohsG6T3hXkLOLMZlh9ey7ya7U5P63cq046GDcKUfZ9sD0BNSNYRm4rwgZJG
zgI1DtgJZzac/LJ7g7kUK25NY/y0Jwrkn856Kz1Q+OfmU6lnqt/J/p1isFBIHHPW/UrMcCQ2zNM6
4fVJe+KRGKc/eS0M5kNm09d+cElRKaVKqD3ktNqxz54R6K3EjsQVKaY3tHa9EecrDwI0KUSB2gWp
g7Yj/vq0AyZZUEOsc6+Efo4abyHEUJtMJ39T3zN+WN0ng5mHYT/k+wdN9WqL0CBloLQzNFJuKdyX
AwwD7i9hq52VQ0fM8/yp/8a77BcMMaeZ/LiqYY1TmqjG74nyIXvlbF9fttT+goPToVAq9yFL0WTK
e/Ta0sbVgHXIeEQa1g0q5+FhsvEvleSTJd4eyOlayBO+Xx/UtbgtCwpqAtnxvZ/gMEwiT1kdcl4j
SEUXQ2Kpp2JJZDE6/B8SPbKsf4iWu3XKmBA9rOSl0M3InlF3FerEZ88vLMQ6UiXna0ZRJQBBgojl
qrWLTnYIkX8jau5fK3XcSJlAD7ABPfON0dZHebqdWrsd3dcn//1RPgdWf3Qfy0Fv6jWrY2dIjx1O
YRpVnyfW70mGth9R9wkkWLJ8oXFPQqWsP6VuqgkF/kecNk++dvZA+fvdeVMHlVIurifyEnmMIJYh
gMjZI4GTPrMlBO4ZqbnhvDF0eI+RnLbr2TRkol96F/sXmVpX0MzhZG4b2+12wEdIEAlsUehbzvpj
ls0YmB8QSkTIaEqCqmJfHKo2Ti+5Sx+mbqJhqaoAlx4q6UN57+Om5pg5PNaI+tSU6FE2lG3olshs
EN8vBaZpvZZT3NYe6SJ6Ng1ESanws0BP7o3YAY9WsieG7CIKdgnwcGlqrR4O2PjSD1VJVErdVpuc
b3H9CTHf7LZnqnM3yBIs0+12rG0LGp24oTAhptBi4sRh1ERo74adcaQ6wKJXJP3KN3YpXasaqJpc
aOXQd+C0bt86jxmYNtUj+JTuKuz0oZ7vZnepHwhLgcvlwXv1wPVhAlpjV0aPSaj5T0F6hvqJ5XnG
uAZW82KwsbqJKo6mrKGYnihAHuJAmHi2kQa/84ZMtui49Q8VYDlsI+TeruM3v9WwAvaPdnzJiDjz
QyCTCttwQ6q59w4CSVCJXCEob/y/GbTE3tGO+iKd4Y3MHZAbqXC0elThAFml83jCaZY7EqbQ/9Lw
FQiSGiHZehsAMklnlUVTZWwrlwuMzbaL6B2A6dT05pBRqbg7GuM6rY6DVgjpago3YYrfsboUPXeo
ZvJ2u7HVb/0ni3o1kBO2gzF1OVjLN4cvyG++e4gv1g+nxWW04nppmCtuJ43N37wm0dSKIiI4O3nE
azLKeB+rqkMhoK/vxrITGBGqN22c7p5KjJpNspsIWWnUAsPotHsvBKwMaKckCrCuluEYLLYqgGJw
FRfYMweBq782fbJ7CPQE9zs7ln/c5Igi7IP3i9JMfX/s0qHOYmtCCYUnlQDhXubZ8MlRjXx++SHH
lDpHR+Of7DV8AX0VhCj2Sq8M4lcnEeT8ljcS20l3cV45Vu6ISSCr+JHqJd2xCNQyFKABH3VGngkO
kOgJChk6mwz+ULsi1AGcgM4/56gW6DGo/du+6cL46/bvnYGQjACezoDIzfkH7DawHvMbfDXnIO0c
wrnb51yE28yd83b6xmGk+nGcsQJcy9oGr5/mPVaxqLe4a7njE3mVfxDlKEY4pylRx11OTfsuDhWO
mwVyzSIjlp7Jfg9mJkWBCi5MbaZoLAT6d3E/X6CGSp07JYDi0YrR8ffud5QtodNj5/Iw92sPGWRT
Q6D8wixvZ3zm5YCecv0QDDxXoTtSHOeqNjQeOlUopm4dxaJnh7VZ9f9tevWOVrxb6BdBUpJ/dzBz
LtevKWdSeh5lsdM3LWdY/FHcqVv8rLsUZwyvMLZjRIvcKaqP3RDQYUy9Xsjay086MVZwYpVUJia/
9YdGRGaEn4oY/yix9sHlVMg8oLNgW8i6fw9xKk/CdgUvPu8Z//7aYEZQv0Yk483ILC58rlpAh7vd
RAOMK+7Il4laimxGuV10EaGYeZ7TQBrvfKmV06/ogIAmaRpPW3EUosBAF96du+YtpcDP9i8NQGq8
iyy5y+qMNTI/h9qg7vfxDxsmeJiR+et/LOrsZQcxGh7Ovlj9x9q2LG66d8mytQgyMnjDeTwA259U
qUjHjFYzLWuyiZ0Ub2efybbRcNgvw3B2ucoAnK7ewjZjj20B+91Gnz6iVkSldqsskheOhPIp6f2+
l2Lg3t4NL4RD/9S63b+qx9sMjHeYsVzvIf0aqsLOxmhZY+SFdLY/6VTqci/BTVnz0n6O7MK3Rtwi
yPSjfi1cwl0Y9dY6Cw8BTKokYEtInA2YPaKcegcHtgnOthYBYqj9A+GvsK+vMDvoGnhKFVaR9kyf
JW71RrYp55jNoQNf+Sha8jVyEb0VL8wM6PRZmJiiZxpjUAig/0GKXnIduJvObEzE8bbyjj1EXtf4
CDhh8cTCCac5bxZUIoKmI+RiSHtxnYOpkkS6D8wWKlJr07p6GjowhqAtyHloCkxojG9/bK9v/0yM
wK4b8RHxjAJVlv3JTUE+A35YOrUOMRTuHgUZYUTyPjNGXc2n9RvtlhhbVhDDbnU6XEL+KASt9GiG
gdW5PNz+xvxdStHMXioH6FIgKwbJEuqTbI7aOOarZABIVx0GNZgvzo53yXplD5ALoMwg2Rld7pAs
/TNPrsqjlqke6qpC7vQ/NwsIL67Wv2UpEvF+9kyXL5lGtQ2tW3ObS6mWSdQmN2gfzaWB8nfW3txN
oDJdswn0UDN+9VlLVTPcRVgvoMjYVS1eKWLAz9JSYiemeHmh8Z1vZc3s+Uq/6+TMBdf73IJzvw35
f9BVO10Fkta5e3N7Pn4PXUvtPLkr072lKx2fxi4Uqarr+kheV2TJuXGv5nJuwo5ZAG2dPqhUVbND
3MWjjVz0xdLmTQUagaTfNv0APoWlBHDC3EycpnAK3iqViAQyZ0bzXe/D2i2bpRyRPbrbkvbvTuv3
a31ZlP4HoD7hFjbtSq2N32ahnpp2aJ9bwb8JTTKWfvXucVc5VXCJkyJVTeVCLl5YLLyD3lhxXGPi
jny1xZGC54ZturDt1al2GRXE9iIbR8c6G8FHHIbBpP9l/yixi4oYBwpSP8W1kr2Rl0Ime8BA+SH1
/gnqLynTbXtMIvg9J1sG1y1zadVONsLb8gzS9xw0hcM6mdtbRkNFGzrV1LnVGE9LXpUYNGeJ1agY
TM75mtWPoHq6KfYYpgEEjyy6wTz9gG3pquGDfk2Cu8KDs3C9idLDwVDceLQ7etehdv++H036kGJk
HJNMtmrJ6NxzfQCVoTzjh98QmQq343FjeG3va542jwJLlTP0ftDmhtqsJoYZxTpr7qqBKCiDIOrr
9PILqhi0VokMSGFqEh3k4HNYGx3eCB3eNNYZDkQg6xZu2+aTthOoCdNeTYrChiaRSuTNCgCRdXbK
+x4PdPObZ33FxdVHIKL9Apwf5RHJTZdVUpIzb7qABIxy9zDQ6BrAbu10n+kKS1534TV8YgMvYLGF
E9wRbKiRDUjl8pLPpuXNNS9vd+cuBeP49z3Ap+s3ze9aL7ADy/0/pwB/X+NeppMnSD/ynLzMVtgw
ipu13vLKk07oETwP6VLH+qDAv4ccRQQpjxjWGhHKt7j8svD9YFZYwS4EsQ4g4SWKG+Bm/JdLE9Gc
AEv9Bwkt7tqp7xSC3pZaVO/1ZTK5AOyaIgvYX/v+5GkIsJE653pWMbI6tELtfQq5efZKtC37NK9r
l3W9tbMhrS/oorPbkbtoX3KuMj2z+5lTSNJ4cirwvOnjqVs4S2GWMgPoGwj7wE8kIR5ROMPiON3T
UMaUU688ZKKF3w/NlVXT6ZI7jW7s6WUTSbua/9+sRvC2gUkoo/f6UWodkP7+F2kR8k06QB45Kvjl
rB+Lim6WSzG3Twi/pfBjgcIHJQUA6RoHGjt+JEf+Uyp0BKmMLGZuJiA28KZkOjzanMNyz0Ibb4Y4
O6hfxgGckBPZ3WnJhrYkPseM/bKIqk3ZklaM5RW/fg0cNcL4KBGLi0JGXp/EudC5SVih49cZ+DWc
XhDQEh9ddRU9LdXxWZ82OzdEIZjVR/WHS82FT6oCN63NEX9AuI+OlU1835jrjq3QC15Hp4mTaKyS
Nmbu1ALRetvmnBgKVEwYTl73OgroFBrvLjBlredigVwpuB9pcTtl8I26txvDxl7DlD8HoHoyPaZ0
YIn0puC5naTbMcsv55bh8WWPoF1ASucEchFQLid6LOZSfDxLlJV7ASzsVAq6K90SUtZqHpWurkGL
Gx9Afrpy6tmyz3zI7Io+Sp6L7xi0YfPmsV9nH9rlSGp+j1ZohMAWpcCXxgUg4J76kcL4IJFPzkYS
LtVk2MQtKuurEYe/jd7bTBwmHaUyl7DZhOoNPHh06rrO3/h3xJxPifhMAMI+uVoBqKUwz6ngYE+A
S+g3JLZ68xeiezL1Q6+s+xkpRoGtMXgD+xnRIcJdzf2HipFwg0eLR6VtaCOxEpOztWUdy7v5i8n/
E/FvLQ7kAOagXasXRf9BE/haL+2+mGaDOCrLr0m+NqhmDuhsNZ3E8xmE0IHapPOKdm8ZmQMrtyoV
ZFVnusiixRv8PMNRXHm8w5Mx/xxsZGiq30Fv85UC5u7a6XcY6VpAuWdGvmPkZ6RKKOfUQolY7rNR
9upU9e8sO6uj7HFxPqelyxPCaf4o1jKd4PkcH+l+GhqmyhgeeRCGKPSPf6bgrOjFMJnWD1J31lsK
JUPzFJuUE5pPaFU4UO82DaRWcyFaiH7T4FcPdyiTtXbOIP/s3yEyyxtQW/sVzq53kh3/wrphUOnM
3zHMaRtFXhoi0TB/L2jDQaZFxqxOvRruNIukdI6cWSrVhEl0mnF21ARNMnXcWlrGqC97Ym4ufo0l
zanr74SBuuXGvZv0bqag2uJmTvYlfKRMq2CUvysNXTn/qBhB0AQnpS1as5gdGflrCyOALEPhzePn
85afSi8LQcwnCMGvK4mxgI73VQ2P7RdPeah7eG7nxVKpWM+AMBOJ0Sovjw2AiMpbGkefJi51vJrc
rjkcTN7fYxFXOuhw7+Nq3CcCLfcEWeWXBKdPr4oSDnH2G1lqZci9Nb8ZuIQDiMpCUZIW7q6F65Ti
fpLlm4Uhk0miiKHHGJs9iX6pX2O2hjGrSNSzw1ZXLfJNaCD/p6nxpkoXcYMu5Y72qGa5t4u1456G
CgKjDiB5arsD0bccnUVGh85a9fhjNPA+3w+Ofqy9ZG+qISWskIKm09ane1xeUarnLZSb3CjpaZym
jUYNdvYW4AHn1cY13DzaOpFRbITb4KpSx740a4D03FjtmrxxFffqA2kDLgU236EAwHsw8mzF/4Ub
Cz8NVNTcPnKi1ZZl6c7Lj05ZVaWpOYxXiM1t08Zds08BeqWy3GrISsAfPV/9Nhl81MwCZfuqoais
t+yM2y6c6Z3Gjvzup5SyeEqShBvL0PNagiQrJrFl+gJdV6Dcs6pbU5gVCqbm7ZuZUjQdU6kaJNhD
xPgpYtmz0h+mnj3gdEiNwWQb1IcrOYDIbmpiCOP9AJFskEql2YtPt76N5ROOqweNLfykHPd7df/G
B/J96Bu57wp5EioKGAGdN/gYgnSHsRBePV2o1yElDt5cMYSq9qLjNpho5Vjffl9UuPCVBorwXvlF
jRAF19wDf4T2n7tPJcUd4Z24T9mC1iAlfWIdkW1OZ6T3Kh3F+laP8clW76Kz9qrAF1STlAkCxNtC
b4GD8tsiOXyhtNc3Slcrb7T0ud3/CCX4YcHwYsSDfINqLVMonpMN++tktLSiB+Np4pO4AyMLTW5L
4Ph/Nj3yszcyxTZQ72Gm0rZxY2EIXTPKsN5weyb+tfzvOr0bv7frIpQMA5qvD65mXyXa5LOKBFse
5MTFLebRR7yQ6JT4T4le24vcoiHxQ2x/4bOgxoNW+uwxclSKLhFuWisOvga8+5/dd5vwSXGTkAkI
exJlMjDyPB0Ms9iL+l1Qn1NebYnVWEZmp7/9dW2XgsrkKdnzU8SMdu6jDjA0xJYlXKVerjDRaZFP
MvzJif6UIjEEMWkb6PTVqR2XpHSyIXKuAd91F6v4VSAl+hQaWzZuXSVtQxPfGIv6Wptle+bEpxDf
n5qeQyw14PIJFQmwHI6rNDUHrCqHO/oE5g4pN1Cfc2JUY+eLiJuPZ4F0E7wn0Av/9gK4aF3YxuSB
FVfaDPw/RSwaAEy1FjEwluYH3IU3KhvgHxBZT2Px1X0irmJXVavH71Tf2CqcyAu5yzUFs1/99KAQ
phwJsVCFc/UImGOIrqtxsHRcCaS8UZPAy6v+0dw4RMpNj60Bl/bh5fMXtc3brHBtWC+TMsp/3XQO
nU2CaBrs1DxILbPr6o5axcZmBTA2V6cFKyfBUJJ00hPNfqjsP5ENoqGf9fu9oiGtlZGUEeR4xDRb
ALriQAWtFNYeScVmPSolfBQmmm9MIG4gBGFdjWz2ihrJj2Y0mC5AsGLyhi50ehKySL4Q+P4wA4l9
LbV5AGaODJmWq3FJSvV1BISdV1u7flV+89sb/g1hDqJRBHYuYcsQlMh5CHNaaflMAlqzml1iW6ok
WCHQ1MU9YgSC9vrMi3JwWDCCuLi7tGInSBF9zZ7PM3QE4yRGWv0LRUkCni/6F/t98ttF4KKBDkZa
yP3uhpVPRS9sKz+riFLeSajxSPmG1arfbOFIGONLM72pRfb6CKlPSX7dMB/pXHc6px/MwF6YYXTC
zg0JDk8Gfp/GwtUhlP9DGWIlpbzG30R1wy6+Le91BusQQBey8Z5vbGfkxITrvkU04hmazq6ikt25
ZypJ9pMWeiPrmvHJu2WBSL6AeUurM0SUN/xtx5pdELV/FmIex1ngbPMpoi1CYfppI/viRVgZklkz
zgOCQJMn6V7T4Pp04Tc3PRxnFEP69guJUiOALOYj0HqBYDiKqgmfcVGZFKlShCYbdbW8T7ypmuQZ
ktpFpeQ2f6xLiWC2UIeXQxc+9kcbjyZf8CRtUpoJjOcwVqjVJGbhmrLdQWrxtYKs3mwn3OvdwxA1
gXTE1BUUwwBMh0qSb3QB5etJcph+enEWi8Y3QBD7h8OwX667XScKPCZm9cmnDw+C6XKjTzAcaTqU
Vma65Mc2/sZvtWFWJ79+KcAV9FbepaW2WHEOOT/vN02IDX57xbRfC5jqwonDyPUWs7njj8J+NKCq
K1nM1hLnkrbIyd2pl5ToIsLKPFrC6VBNdQ45wyNdt/5eOZuaR41WFVJhbxN4Y/54SnmtFM9YDqSP
V9BcRrJoMJ+EluHEhSSydzxw40uQfCYYd9n/GsYUeJl42Y6szeSgxx7n6DDvjQCaIGZcJFAgO5Ec
qh+iB8P2HADewMs5jzJStKR9jrwDnvnFFPF7UTMWApuxS6vzWX2utoCO9Nxz9V5JvrIUZqALVHVo
9OsZNX/QVLaB5rOc304hG56TcDGPV8W3ax0AAeKZWKxs2H1Eaj2AC3X0cLXVMIdf/Og+I3Pgs/zz
LDdKMiP9CDQNTY5B9aGMknTM7YE/F6iGXZMIbSidFGmcgG/3KQXHcvkESsA6ABJA42j7EcIZgAon
ROE7s5LQryWbWfL8lcjBs1xuvGuT5REDDf+FKYZro1MwaE+FlizpVErB8MqAdghMqys8FFwUGJn5
d2Eq8sncxIUBH2JYuy9nxApAjxu2zw9wGsn0JLtfUFc2g6vAwe9kzbE8dzb54ZbPFUGiNICDfOUH
I7IKwGwGZgLuEcsTibHOrrDIXTZ4n/IiYWpmFJvbD481T2L8hDAJTRltbRz7P8gzyP8tuEKnhpiY
mijaHUkWK0PzE5QUvYu91pEIdpcGntViSxWAAlXXLjSca9y3OCH317nieDZobo6U79IZv4j4NGWD
DShUMJnvNd9i67l6pGOQDOd3N0StsEX9e8na/ox90Zcv5wpbdlekFngWU1HVrHD4o42HodymFouX
g81op/xvlFXb0rIyuPgsL3QlGfXGMfyc0ZT598GOKJS0VWd6ocw/xWPKX5EEndpA3tl6w8D73irN
hohRsN/tKKm/UZWUkNNnBlcu4Q75IRfhswpkgmG8WYhLBmjuoOr0jsDE/hww5fVS52EStcKnZAnK
iXAuG1upK/BkKJuV+UdspR4a5C4Z1UcT8e1CCrcbp6Qa4ee9NCjJ/S8MNBHXWdEypxYQcanqo9iu
ALHkYwzFlpuBplPdpJwYK0PFI0kBDIflm7WEIgMeWqk4SDqwIqrBcLqN9xX3cvp0YD+MO9+aEdNY
7zz8OwDTYe4VxD9MxQoRBKMaiQZ8l6iYiVQSuncd+bbO2rJX2qmLCwJi0abMhQWskX8hDa6yH87J
S8/V9U6NdIu1uNubeGkj60JqltNPsOVIIQWN7x6Gmq06Hax3B+3MBSmk/7X2Qaq1c0qZIczEPSiJ
cHnYaBaxYS2DBd8ouiTr1xmKBF3gne60etRnGG8a9+LnjnlV2lt9Cio2b6LD5nnL2tnfT2+gmyPn
whVLF8I41Dzn5FeYrkbSPXMhQ/ps6ILqAKSMFenRzAVUOIwIAJne+1QrU/0CL8GB3AFvrcsCgh+L
RkNViZ+2q+Anr71v7Xr3+R3LxehdV9eLOpqHz5SNTb4ll0dypqHTJXGq3QXFIdTTPzVZvwYOXejN
+R7tQn6PO0nDVDvsv/XXAzwK1IwPvJh7TW/VQ6m84oCuS/+Av64+6mRCtpKyOevxO6QNvcSCn6hX
dl/HHSjsChNJjFJ7Zlvr4IjzLpC1rCnRkGFHYHKPjuPv+FeZ7T9lloHe+Zy/FdH6eCDghvQFvFoY
idS2UUnfoauxw0AfYxhoRkeYAbsC0QTRdnYqWkIA9wUAvKU+jz4ryWO4E18csKqYChGkYoC6iNpb
Clt0ZN7JgRqKYUz+DYp/tY0ntHJ9tZKn29xJ5D/bQB/m2aAA51I+URCle/nYeicjKNUhxJQfguvb
Z4muxqGKJ44Vkx+OgIwhiSYp9JmgEZx6M2qYAvFtEr9R+Jix3pyzJ1VOgic17UZTaKwj3PNbmz7c
HN38ZaJemTfMlzikWS4SpDFnbSI/Y5/3M9gG1mOg4s7bz05iWQ7LtiTEyUafZfD9/wle5GfOM3HH
CL+RYrSEZDPAGU6Nl26kiAdUaGmpsLszzqDGH2y7P6PoNFAi4D7wuWeS58rBZ9V6eV9NkbqLx+uF
HqNJSC4Z/Oty+yzeslTl/fKnwgrvfzt4CkG2mAze6qt00B4hEIgBpwcOFRq4WnQ+7HIW7y93XGB/
hOAyeImXZzBW0uuPWLJlYaMmZenXkWGEFC3SDeUkKWRayiralLVQfThqDI5ZGSvFHRO8zQN0Kh/0
8OH53uvdFEttLOovk6KuTgecS6XU+1a/TICBBIQs0Ms0ceDaHJvQyeie4rEqjPHKZI1l2gGfLO5i
XxV+6ECg5JFl2bLI1pZVd7kseWDKB43SXA7buRhTEMeMEFTMTafi5QPbIeq8CU5vLH/TS2eh0Ny7
mLfvz5a2KbtYlciHqx8RLKpD77LOerMUdJhggvFaH82OxqoZg6PiGIFHrm2Y7iiP1DpPGCiHUKSV
kxb2eCinhUgVc83bFfej2tk9HN19MUrW0wmaAbta/kBTUdWGJC2i/XIeBFV0dkPcN1GGAS8fLCxs
U4HB6t+Fwn1uxEnzbE6j79OHwjpaNzuRGs8IBLELynkqyKGdr7188S7wIDYGpz1RktiDBy6lMSel
v3F33qFeuG/hzXd9jFaM24tA39u3ZQoGXFFgmTVmnKS7i6BwcmQWl0uAQHxKFyQ/3PxuXUK6QO9+
UNRqs55dPcK3XJXR0k+4y+NnC+WNdDJnaOEf5egPMgC/DpNFRh6rSgS0qPgIk1qKkwgwTB0/T+F/
jWDKackqsKXN2x4WqPsg/Fq/NNQrOlx6LE280xl5rXi2nJVnP0WHfuSQSpQxtc4Uk3NxRHX7n8f6
xSX5pF/q4LZVl6vQ1OemVb24HAYrGSBD/N949Wv9keoGTU1bb6ZRr9oY6iTCwJwcyoPX8/RSe64f
P19EZRGeEU0+JNWva2srjcSR900wqYeiGy1u8vNgi+VYQK/BrGXW2vNZsW5SrH6z2hiTy748djIi
o9iNyDEBaJlrliCKeDHua2uHAihyDOmA33/f0loDdtHbJh6LCUINVpdfkpVL3q79/C69asj3XJq0
jMQ/wwsoICNYrm6pciuW5velBtG+xh/4bKAMjNswXVwXlCYABeiSKOnCNPdyosxWU90oHVJikf9R
pq6jzMRKA60dfMPSWclckTIn0o0GVzpl++irpxQ71sbsadFefdAghNTgsYxE68ibn5mjQ3mUmPng
O/xy7SqeLhR4K45Lcuwp+popIYQXfsPECNlbyWLjD9Tai9PM7PLrLrApaHcV7KJUhcqmzC1Hqop+
tx6iuE6kdNYkclVtAwc+A+8GJ+aDy2C6PAIMPB4D9M20rnqCndwdYLXxyDj381LVvOcnVRYBFdhO
Mb/6t81RjzSE9zk7O0HiC+daSTJff9M0z9oY1Vj72zQcMnFxH+xirrHQinbHflSNi2kwbayeEx2p
xui4Jlfy0WiaMiWIqFrzstj0EF47AoKwckw3dZCkcAGmjsAAZjs3i/haEfVlJDT+TXL+S2wAbTi3
mdJAGQRlPjrUIje2RwuDmMR50as20dAEUl+ariY4yLXTA6sFx7SsIcCABhgoiz0EZFCdMXyfXjIO
M+iaGm6Z4BgLYytSuP0vUuoYrfF7S1HIozKFHdrfgot2aP5lUxg+OLFt94HMNMKrSUbCkmeAI4/J
WYWWsGx/17Nm7IjA5HZggunE01cUrIrZa9bqtspYQyptvoxIk+WPvRgO4eqcys7XvvqEyHEAfzUU
0Dave3v/qlxOQG+ds2lIcIJu/q1d+/YWwI9CNYKpfQPYZ/l+nKJ5CwMDFd9QAL/s4irLBfUaTS77
jcaEeHO82XmkoglLSN9S5DpO464F+e+rALoz9n9a8yhIW4WyzT+5hxRmGACpAOyN62okpFLMFKHc
TwY6+Jc5Kt+4c/lfs4EfgnglNjIt9mHrOIs5ZVdtOsbpqhsWcnhwynlQ9STe7YZM9Ht9LbR2ENIk
nPpVQRT+HrIiYz4bGb71tgVgj/5MI8nXOsWTFtj97ZBZCRqZ3umD+bxRtz469IkcJykAh3veaDEC
hP5/HlaxZ8UNY1pRIdTE675h1CceLpUQ8ABRBsnhmthF14Bw15zqsldMpOXsTdUczrzrdYjd/JmR
/5H0tnlgHzqZfivsXkFbgQnha8tf6lsADgxpapp+RREUnbZ62n750zgnCvT4xH/UWWWIBqhdS7Ti
Aw3fWhV8xBCdTmSbx7/RI1kMdoTmgZRMOlzBN+oAl6tCd4QJ9kz69NhyAQ72wpfli+Loe/h8yJl4
u0iJN0Pm+UxyQqKBZBSkAlRd37h+FWxBJlQsm/dpDIr2hd7ZhBbU92zwomgFnibJlrrFtJXZGpGk
mdtkVOXvfDl2hvZ+hLDYHtKvTwss7RgKaFPJt+qSfJA0aQonv1034KjtaxjM1stPkOq/UaZlfRQ5
gtHU3GOQJikaMOclXWXtc3F9ZH2U4gTzDluDNGLA90t0PZ0IWIYV14BEwyg7L3kbcfUKgXUvqZ+R
oloxCHpubuXUXiWWAxZa4aF4AL9CWJX06azrJDcdFMi9dPVwW39iyunm3XIv79BlxDSeczPPpFsU
qec+JjB3En+VysaWSE9V02VaV+Yy/Iq6oZGOjgYe7gnWk29++ffV2b6qOsS5BVZiR0RLvgzEg++q
aOZRRi2PgWj6BSgDlFBXiI7GClkL9rSH5AaxqPCbLEKNumQ138NzoMmsQqALARVds6aLVlE4mL3b
KN1/zjCadjfGba9WzvwNbzV3iKYyBjRGC7GDsUsdBIQf3NTDiWJ/73TU8j1hHO96mPw+vnIxUYqZ
qQ3HF8ST7GujN/fYbcZQHovUnMVmVegey82G4yg5TcMKeHGsU72K+7N0MCD/bBGwxP48dm80+FAV
fxx9bzdSPf+vrd9kW/GuiVWof0VpzhAzHA71uUm53p9YTZA6zJBd4SrwpMx3WiJ4x5nHp1UV5JXg
/+p6ngQKjdqzPXY/2HbmGI9sBaDUXQghb0jzW/9c2SpyRuZErZmbktTCmgR6iihnO1Q3RWyJ/qLq
p1cXd+J71RZ6SAgi6cQL1jSt489gA9NfWH7FzqkkXwrCmm1R9J3kOvo68QKYyNhIUwmVwCQkbBg/
p0Iqey+woUIOHagI4NYfrTNg0ZDcEF3RoNvhbjuZ0Ou3ENxMbTZDzkyp+RlG7IQu2Y3NIjk7bm3o
j6MB5GwOcdWyK3EF84YHyNhpMByLwVt/mV+om/ddOG0Rb/X3gZilGm65vJ8AWMwKkaYIui6iJwjF
4eeKZXXMcZOvG/XDkQrdx1rVwl5pR5bRqLK5JKQ0CuyUAWEeS5Z4w9duiX+35lla03fftJ/1pYwL
QVyy0yzOC8fn4XRsS0+sI5R0tP+zey9Q1wcxSY+YVaf3TU6Fjz3wQo6aVglNy3i1ceb/gWccEU/L
fJKsuY6/tyRLOQBbgGcakLLUWNUetT/ijJwTfdQ0SKYdgVOgnQLkgwyOiSwG5xJ1w0czSpBCq2ig
w8j/Bh7HbdktVd8AR+Y9boosqy+ZHVZm1JGeI7IG8h5OO1uEazgJ8wMgqw9MijQtHmEbS3srn5nQ
t9pChKJLcMLkSnWi7rGrQAslOW3trplsasf1s05seLgVdf5qpZr0BdmzObXU7kkjZlXrnMthm9Am
/lCF9BlTibeEiHMjKBeQZGPhfGe3NRv2/Zo+XJp1yef+t0TZZsQHvrMP+eAhbTZjVZM89QxzTaDl
saAy7Mh2v2eOunR12WuB4zTqeUQBfF38s0QYQ13AraJ5Crw61SFSE2F/DFlYXuiWTt/FzGMP2m1K
iX/HrSmTn2UlLwPFz9s0qeFbn+J1NXXse4bXRjcFo6uyK2xAfWwCbLSw1xdRExkq8F1Dhn+B+6k5
OtIpRwGm0gm5HQIU0JRWFv34clBdGdqHcDpeDNQH2JUkcfFBdsxubIwyP/PGr34GJt9uS6RIaJxc
vECHZHSbOiD0wWE0DVm+DqxghFIsvFHJPaiFej4zxD/OOsuwNxT2lF9JIRofKN7CAmL0TH5A8n+h
EW6hf6dLYoaBbSzdHI+HZ7tXDhxht7x5nbqDlfv56w6wDUZC+vqz15VVZJRzt5v4mKk6GUdcCSA6
3c8nnVvKUw8gFU9kmdHf1q9oNYSv4r0tjljjjVoZUYkGG9M2u0c0IPyLwusU1tCwjEofGxOLbcge
8cOZ5IM4/TTYw11XVTwU/G3Fi7XxM4xV+CKvm3GLCoBB5iOv7xx435tgMB8r5vdH6bugOOV+DeDA
YKUd6eAZBZNBw4t//0vJZpwfiqcXc0JA1EpDNAR70GZU5/f9xqgDLA/TFCOBLVEY9wUd02/784bA
HQ/O+eOI6RGbCz8c0QS1VqK89O1JM8j0SEIEyTm8ZWqmRvyyqR47Tg8X0q2O3te8rCdJxtC8dFSx
5mn4wpdBQntKlB/ZFtO8gqbCpE4ZTE8VWI5Gr5K816aI0cn7jH1KmAUO+LvVO4IGel2BY+uMRqk2
6sou9NImoY2NqNzNwO2sAVmVWFXH3Y+3U4SkZrqvoKXTb79MenWnA1AvjPkI1DWBhoKyaskLnsF7
7V+SW/nIdp24we2hJUtZBInNgcBYtOywKLAG9tUnUtTdcxPHAVif93RigNKTbR5IB87soRJgQqKc
xaj98cfPE5SQu10s56J1n986yOdL1M/Dan7Sz1xHg9M8oK8qeIaxN3LdVhHBZuw4fDZ8ZnLIZ6kY
vdQ6ala/w5jRp5VtcADhARFzl0c7LDYd2iA+tN4KL9miPiIZrQs9CA+m7SnAMub4hIMJKfcH8vBY
xY7BSCfCnW3U+23+gIJ4X4qkBbKX81bRhAADZiX6A2QlrhzJQofDRbaWDzvdKtI4ElGLarE/DLk7
cBz/z9U5GvAyJO4qeYCLkCXOikfUcyGvEIihalc7vfL1zcFUfNP/dC/+bEWC/9onNfl3a4gDPC+5
2UrooJo1SRyS4EkHvDENU6IbNDByk4OMA5LrFp4fl9dLImMcpGtf6XVpbNpqVOqj5xpFXk3CqJ5W
al7/p7lbUzblT5iZPzYJbsM5BS3Xg5WyaAroJLD7iqJKd+2CtqZ2XLgrm1Lf/6JYem2pz0b9mcCt
wghT5TkgNB9INL5FdERUHCUHpns9zrAxTtrgvE9k/jRHTwbtNfYC7k7079Iyj1QRFTp9JzpJk976
lEDOLoqJnAqbKUK4nBD4XhW3JlzHtaXZ3SnMtIQyDSw4PdMSdfTAqVyvIx2EB2IUfrUC70odCv2I
13cM7l9edKZsR2tBg/n3WXrnaeGLMi7hy0ih08YCZr/pM9wfnrf0LyIPJwqTNlJDOcTxFsE+/CFf
hLgR5ctf7BkgDxQ62Y4FCWrmNkaAVKD+hBWfHuM3WReW1iuuhk4NbK0MP7CUZ/LDtsKtuMnE7MMB
ulqA2BhywpgwRLAIoX1eIafbp/r+NGgldCKUd+JNvmcUjr+c4mA1wvSPZf7Mopyhjqt9saQRuUk5
HSUsNF6jyCCtUzOQFEeJH4QeaFMPbM1kWjuV/Trfzr9xeyiYo1RKXAXmzC94W/AcO6lGYu3n0/Y3
YlZWFCq5uC9kSsFZ/CxjEKlRn1dtqoBYqY1UQEE6FAaMrT1uRuYJ3jCCJzVHdoDTDR8YOVXuCrL4
0g/YxkbWp8CLyT/JkJfFZxX7iXP3wcQIGqw30qKYMVcgAyc0SQrvctbniKbC0esXZ9dDFS2hxE8Z
GdQZ06C0GShF1hr0ri0Kvl/uVCavcxkiFqUWmt6wTKwXVP9fBDpALj5aJ/pbalubVjMvBJ7prpX2
Kkd9fivvTeA91LFYLQ8aqbp5HQ08Y+ybiBEp3EFm43HEE++3as2XGCkHNZqUKAMyUh5sJyPnlz7D
9J7YmsUAXh+DMxK3NN3DSZB9/naVKhF8oEbBBtTPJ8ALzc1XJevcrRsNBTVfPgOaDpHE/O4Z/QjO
qHdPB+s1pYvRrVGPGO568DlKH0Ys+M3Kon2XZiQwKOrO4n3GBUei7YIFILDDZ8A8kGtGX9+JO3WM
iGhkaVPFxry1wAYOSW0pbvudvvk5QpbhxeSRiRBWjVbyjp0NCGzcP6MRYNil8B2F1aN7gJ8Lho7p
EO4TZxr1pL4C1cRhDywSD2puzww5lRow9C77U1zUgw7xIFiWhy1JC9NqERVyr8IYnsp7gQ220Z2a
erStDmQc0DqnJ2/gWJ5DQc+vtneTshIwkx+AEQElePoCGRIP49e9WexjASN1bDMkGn/LCxDS6XwD
+LcHBt4j0Vqjy/9YmoZeESUd8Zv9mdnXLH+Aw2m0EoQFRFEk+uEXYpMkNeZhChSlKBSa8AroSvbD
C+FiaWEk7oYQ9HcQxvq60ogE6Vu14/lS6cFBp9oUs+q35wwiZ9SjZ5yy0b8HX+c3SH/3uP+4l8Cc
rE7jgavzJFpPbrVlWPub6pihskpE6MM0XrN57LVm8g5jZ/brspRjvUUKzkniXoCORnC7n54/3BOf
FdNYuXoxw3sOC5SDAo4Ub6ixSrmXhnCtSKhKDXnjv5Flusl8tsK+GGlNwt6ySJdS3KmKYsr8qjYA
2dPTrG92HPmDRlEwescA9Rcpvjmsy+3NTDmmu9DASWsNVhYg44qDilYEYTNjyIim2cf4iN620sLe
lgKYd35S1fOq0Zu5q49tb6UwzCJFOqFRYXbuJMcR3YiFU4OFLFEr89KfRYO5fKQhxY9TAeN1tgsM
ZcZTSfrvsLsGIVXCpdwPZvcQPwvRoJH52Pxd4vcVyejfof7i7RCG5oZmvxhE0JKOwQ89NPRAiHgo
2wLeCWKRN6KXZoaR8dNQTXG6d7PEMi5qR+dcwjDQFcDToAcYFuAcaoSfIYNhyB4Oi4zw9UUEvScP
nav0CPOC+rKIZXKKejOynPUUe6vbq1Vvm0TysaxQePkUhiWlCS1grCHdTyKevyB+o5nkXzP6tUlH
uBnV7uNQyJmdk9ilXi1zlhvuJmP34bHnazPyDG6dvh/9cWxSjHeaVOqkv4HG3+nyk90d8L8Vr0BK
rnUoiYjD8fdBFsSJZQ9/etnjk36+4KtEZDY6gerhgboDRUeIpug5uklJFFu9sUJCDC4i2vb09g3q
5GJ3hkDfh9LssfysdkKMpeKd/tTm7AY6C7cj9+dw5DqlQ9krv/za1jjeM7w3/VAUHF9kDbM2zQp4
YsRCLAnDSxboR7mgs+bpSatzeI5m/G6Gu4hYJ9rtNWquAOlkih7kgugJvsdyON6pgDkCDRa2hv4c
TquZL/zcP9QxiMO/acNmSU2tn2BZPNVTLMKzEPGEGOsi/nJUN+NPxb3QIJUy4X8CEdmzymBczY8L
MXeuqKNB5SJmokd9FhZzemmVYQSUlkloAoC+st69slkAiuMDQzD9RwsTw34Kcvz/p7QJnnQq1Ein
xw/nhm2MZE/u2/d153aLQ5z4p9wlTtHdD6PfpLmSdcELG43icbVwNMsZ5dI8JALe4P+y+3FYQQtj
m5SFnRwgvo+AcvdZZY4R0wZMrgJ0ZBeA/s/vMK8ZDeBUO4Wny/p3axSNygY+dfcRAQ9+B5SmAGgX
kZQ1UGWyU+dqaVEK7CZIETwMVIed8u6XXt0nwCeMCFbPvAern0KupBxm0EAB7s6+Q7p2a3jsLNup
DcRy9fJ5SaXjWy8I2YN6hxQZMpgMBCdhIoXsVJ3MrbAbQNmYzMEsW51Yashv2uwSKP1g45xpFR9B
ZDgdEwJC5WLQEoWnW027BLaMoS7e8Eot4Uq89iq2Vn2nox20scoQlXlKWf2cS96L6J6IUYhEdFNh
nZVTnM4zeDCG7k4yf47aa3IicUjf6cyun7Vh9TsSWbPts9bcxc0N2uIlGUh2sy3L8RTRdHxqorRP
P4BI04S4hjZQN3yNEsqtRak7wLXrL+O7kHOZADEpb5pRmHZT9N2aqsjmcbhRBDXV7ebRxr8Xb1Ch
YLVxXxy72Spp5xJLpNSXt+4R+K1mbvU9nMPO0o73lYC1szWTTl0oi1eNoXMXUDDo0EaZoYE6vck3
cn6bcZgXSrf+57TpNUbufdju4olgDyezWa1Tt4l0GScwVng6F0Eryn0yPC+/40KasDUNBCOPZcLG
yzUho0WiORpdT5ys+/JcxLQEeiUGEwoxE1wlJYQPmU9qBejwAkPUckW8zah/6x4U+r4yB/1cjFm9
lErm+LO3/LoJN2rsvHUX/6RniEJo0YTYGM/DIZlX5JY8SgPNM55l1cjo9QeFCs6f4bJfn5vtULxK
FzaQdXskBEmEtmUqvrxWSYPUQOq1kMiAlEZpz7SNki1vh8uuj8GnUBfM3qyO7GtLdYbrUQ3WvkSc
35wizKUFkdYn07pXhIfPf5+lqgDH5hwkz8cV3wjExdi+W01QjDuehaNwsFIXQQM1m3aOol768JlP
e1EsmMqfUiBhzbO8zOUs3ihoyfQ9VT2yJm1PmixcMm27m40fI2SLc0JEgeYMbaTTkzqyuiArcBUT
s0SKJvbpr9PLzG+x76PEnabmGF5yMF7fQS7xUpMpboAHBjswd3CIaReeZD1tE2W99WpW11668yG0
24lzrwcQ92NfoIyEOIgTnA8igp3jwTWLMVMEJKrR+QlyZMmtTGuuVBXAN9Z7HE/gbbS6n4RqH1Ux
0m9y/+IthorexybQ5EAsYQlg2LFa7gYstk1EUGe8tqox3YY+qSScv2+/qwtVJbJkbslrwfzu3TSl
wknbWSdJie+6O9TIqIlEmCsq1CofzjY8d5iJj4r/1p2FTnln1LxvzXx1Ybjhlvw7P4SjFzR5c81w
tJqvyttPq5yO8TG9KZYAVgwYwu6Xw+qF7mbuI6+K7lQmy/10GD7qTxtCwT3/vxS7W+bA/cyHE/ye
Xm9OVRI5LOoNvhoJX4byELldFJF67NdE9Cg563JnK5aJi45JLdkTuEqQrlm+OmHwGr5gQoimbS7V
r/yrFjismxlxGS3KWh6mqkkn/ebgVaiUSmRE47XR/dw31uk6kj6qrXPCOikEAxLABMjbjqG0TPAe
t+/znYeNOtV0ELGniuWzyZoKUVPdC1oQzu8t8wtzXb7DtElHYtx4jDmYaUhSpcsf7j3mqH8MVo7O
ZOsACGui1XcRTB+t+bkbydBvZ5d4w22bWqIFVBlKHm8r+KMx7qhcDsIuXLYLBJSilp1/amQZbPJ0
EvHBt0k07zYmkoujTIYqPlckHUJO0PukT4PEGcdPRCK4+YmD2wApzmOYuQBcDAJ1nzTIiNMxeu94
rLKeWAw+QwGTBcUHKeydc7qpCiZMiXzKHNaUuLMWiRUaJkZEPkNLvgCtoEC5e3zXgC84pc02YqeZ
5QGnyvkxcY83CHNWBT4JdUD5iOS1h19fbo/6fDXf+Hu7qxt0lbacGT2aQxIhuA0MWyAY0ePylCZb
RBzb7qOTO/T4ZWZ1mLoN+uX+TTrtxpjgMIKytsz7/l+wFIOZVDTUve0SzBqh/zsUlbxdf9+g1SUH
ZiP4PtjXCuwtqiKNBsQV0V4ory422bI3TojiAbRCIoEeEIOMxLJ4t4S0iXcrhbM3XgKEyUy4mTlV
1essSxT/YNIVyF/AvVBfX7zr+gIJqY+xo5cARikOWhFBH8hC585lbGchwZzDbhJQaC7BhQcQnf+A
RS2qQgCIi+n9UVOg+Dd1Lp1pKHAYFuC1SR45W/g5ceWfxt+2QFcDBECMrH1YoG7fUtwfU0KqqNvC
/OJn9ItIq2WXOZAX5uug09DhREySuYJPve85ZbcMFVB8XtzxynF+KaoW2ZxG4ZpauPnYH/s61+LV
DIVRcdRzxvUlYV3kgyD62tKo8micQFF6oMwf7Fg4IcxLe2++l+NX2E+uelvimZ28SMzNhGSLt7B4
lLnb+nyLuLEajH7H7nOQzaCNeLZL/LvwGqkl8ukbUf+3mzjB6y21Hc2q6AjKfKvOAO6iWwnSGHpJ
by1m4TheRRlSAifgt5gWMj40geIPBFSBnAGPPoHdsAMcSJpb86uo1Lv8bbiRLoqG/wLg732P/oD1
oN8X6PWAPE5gcwnQ3gAuECNkLI1AohIt64GZW4lypnq+TjOj0SbJayUBFxZnK52FQ22wVhy/FquD
3or7PScR0Mzy/isFqAj0qOk8e7xeVoPUof4o2sXFslqi989YoYKPY5BMDasJe6mCKnXlTbr37KV2
3llRgsCX/QSGAKqvzHcF+3k1bb63/CDv0YuEJxzVy8M9B2tzfheHjDixOrHWrMLETNjeR+7gv4ka
d8/jyn7tvGfcI5OYhzdtQfo9eipI+LN2OguHfu9xEEhSwo6pZ1CqRR/rPP+czHIT5g+hHH3zTMlW
q0WMXT3DNY3R1HllroPWzfpvA0/Na8G8cdVbXlFinesfwyIaJsqMGWARyaa1Pm7e3qNpNMcOPDzZ
SlOWy2Vc/4tfKwCyuKOATHts5/J95vDSNT05G5RGqcfi4nkTEAI5DSJXySCdZVEFVGaqL2kKPRiI
noCTSUTGvNXouV7pAQ40Y43CQyvh9K/hiEyCl++ni2XIZ5kFzuT5895VpKGKrloJcBDENR0IFY7F
9ua6jkcv6EOrFXz2ZsacIg07TJvAexXe+ydnviiJd4+H08LVNej+mgWJQSfrh7Xs6SqOPNftxV7v
T5pWsUOEa6ok29cXg7lxt0PhLiUEVaTbKtCWRP9+zyISqfKA1yDoy4hR5cux4Nwvkz8bJEv/L2vm
lOeloBAUDjUjxul9DL81A+toWDqOMR05QXkYqtokDYIE0aDpYxiQqFgwVXtePcn2TI2ZH7BZ2QAC
Zhw6iva9VEhFOwq4taoJ6SL4Qga2dnp0+erfYpLfyVxRc9iciSe/e197kmEMYVyZ2FNl6TuT5iOU
X+pkHIY+3t33SP+Gu0njEl5YpNUvnfYcWMdPc7eKEMQ7EzQ3P0M1PMG5FPJGrRHCU8RwrW8mgS8Y
8foN4lp31tbjQx5ydqwogvNgO4+k0G864CwjFlPtX6AmGqSaUb2amgCQ8MmoR/v4v9benX56xfrl
nRUsyMbXwXVkpleqTKfI7a4BL4rhJnNo94UInmVToCRmy53df/qDV21amFQ/ZN/Fr/+OFaNxL75L
J4MOL9zK+lXR4wek0lgF45b1vQSccedVPuGbTojCygh+ZcIt++ZirANUZoPFpHrBKEf2Mc6W1ZeL
SO9t3V4RoTQeoqysE6gVSUxr7Fd7mvx78KSLjNPzwkNXfBqFSlOMGSjKP2/JR6nQqf1NKUKySc6E
wXqpacGQz/W8gJ/yj1XVXf2/vI1vCa4JOER9Vf33S98IEqIgEXQwHdwIXPWxtHHzrar+3LRT8XX4
Y+HE4313H4/aEMoh0dMaQlJU/FUJbcFXMCmToa9AGl3QmDwRBbEQnZZTY+/z6pB9AcfzYZd8xIMi
XSnI8NG686yHSdFcAmGuPRbN+VTKyG3abLYqwRa10kEwG+IvKm6FBWoXwwoNW2JfIKh4kutCpmma
IUWGkIt9T/QxjhyLTLKJRFdmd5tLu2I0ndnISJRj9DKTljbYpoEGt80im5rLF21S2k4yng2/upRr
t6MHYGarZ8IK8jGK5FwlXAvP5nrENrpwC0a5vTjNBj+eBy2f8orzhOBgGd06nnxDRTxN0OcZ4dyT
9lG2HgfHyNOnCiOPa5Ox66bScUI3T9AjpR558m9ZEIJeby2e1YhYO25kSmG4y11U3uVi03FIkflM
DcYir/YP51bd2j5HUkcfdeiQYxXW8CTRosobI1u1SdmVWSzV21w92zA5tq2799+zLHLoXnB7L/m2
tABkrtnAGHpjBashAN5cHV+Y69HOcT9T8qlDayl5gb0IKy726EljuiMbcyc98kWvvlJqu0Z/PoL9
itEELMh/N0navX87cqyi2DhwSMIKB6/f7q+I4PK5JSGLMSxgf/E3/g8laCHivZhdX1Z1VHIk//Zf
EqLxFa/o133xILsOpNKYgb8FfqwyOarjjN5iI+xt2kGSTG/Ktl+dQb/G1jD5Glw3t3rkg0xruheB
GSZYh7mMvPec4LeNpnOJ5sZhse3oQL5CpHcVU67m5baDD55j49atlK5GkpsHFJvFTxlb7O7BtPRo
yRsSp5kkjnv+ZaGVUpmX0lkn0y5jfK3YWnwc6vSz/tLG8e5bG8/vUkXCnWV8r92ytTmrqolZL56U
j6XZaghGUTSToVB+jKdi1ohFXoRuEv23/VfSoyv9B+QYSPH580AM/KopyDnf7wB3fl4iVhKBEWa0
ihhrMI7wWcp8AAl5eR7nar1aPeKdyXNyPKYo5IDwDc48HkjdEc4NGQ6HhMBvIL9EQZJijH6Qzarq
uS5tTWvmAaicqiyb6lbnA7XK202y2BWrTkNp5bdLXovOm0BNyA+eiGlj7FkRrl3vSGyYYcsz74yy
MdZ+0Cv0umMLlChiSP7hZf8icoDA91ozFYkTgHGvYL6gcE53Ug4dQehEIrrrHAdGYIVW/186Qfep
H9eiJd94pJAhsG1EP05EdeRBrQsZRVPw0cqXx9AlaVo7l4JA9f0dQ6AAgBVcmCaFWXZVmSETOD3w
86VWBRcqxu2jB60bH1x/BBoxc23/J1bfDymQ96Ky/kO7E5BjPHqcAMIOiUIovgaOP61h7vhr7bvb
ScBdFBiUsnXBdkTop04n9CuPzHhFSH+pAr81k4MbKxnW3HhSDTqRd6o6XsO0z9fGWfEBshhN7/1Y
VJM1bkKp0kz+wo/nzap81QTEu4YXFkmV8/80LlaTuz9jZlKhX0pWqcDnDivnP2kuIrlAgy8guLMo
fXd7SBT3a8JFedq4xLFvkhLb/Mnb5LKe7aFEeFrlPDaJbv+ddNa0DkgQ0WbZDSLEt+DurxZC6EaM
Wn9w/U6MSdgK8R1G5+IiHQQC7hRRk3BCA5Ta1DJ/RHIr6BmaDU0bZoVVGIMZdknsEGfPQ5JEVtDY
dlMl+glzQFsZc5LaIvAkDGwmHQouXECbHzu2cIzxrg9Ug97/2Jp9FdzWGz6ZdsDz5R8bIaycCmLz
IBvrJU1n/yTO5D+drniurmEfXKi+M1dYKdDRDK1B9T1k4BjynlInmhQx1ADsXBNqX9GTJD9bdNu9
Vs34esJ31M2lMoML5CTjQCJEf0KkACE3yWkUX/JS5chIrvKB0Iju8sKxYz5jCwtESc5B3RjRRZ4L
9SMiwJMOyJ6i/extPJbioNE355fF1kqz7n66oZN1lq99y5xceFQuTLLWg7+9LNPKrjgxEg/TJCgH
Ti1YgDj4FoT6Hjymn0jUND1yPphWJ+gYiX+RlcsX0jg+4rSaea5IoFGAIHugmHhgtWb7iVC8qzxO
AvJJJVUOTDCkbFPf/gCpoRK1mcPlDcdRQLctw0kyvpqnLc7cq6UUs+bdELc1vJ3w3KS3vNlZMoY7
Nir2WoIfVR8/9Ibz/eUq3dtj+oAu3nIbjfBXZJ+523T0luh7n6+u7h5Lu7KQ00orhKa39oicXBnE
qR+KJNtCWyIm2eBIl9hOssogDzrVd9dANs38JImWBzIl3lYaNoVHcOtvsOaNd1FICae4ZwgyJ+1Z
YnlhLTz7D5J4QxWBbYiJR1R3iW/1NuCJeGO3fzAnH+HhfZnJK0dJB/W+38mixuDcW20Ste4l/D8T
86eB2Va7s6Az5HxI+fQ03ua9etUjQzxG0cGKwLSOwhi58IEFeMW8vYvOd16ZOl/QPwiG8gZCPcoB
2QuWMgMTvCt6EbcU8Hr553dLNGYknUej04Udv/MX29sa92ZVcT02HhS68s2FAe97j4BJS+7/K4B7
AGg2FoU0rdcQ/oR1stFRWQJAdfzEegMPfFlfX+gMtGsmL1ma1a/+9YCLUBFUXQmyYrRpD2y6DkWc
EDqB73Pkt6klx4Vo8VQ890MuY84hcbseiaZXhtLZDA6ygPE5aNCXpWWygbMAmkSTnv7MNRdNrzbm
/4PiinUNXDSQBTc11DlKIYzqqM+icRJ1shOn2nBPbRbzQoI3GJSaiiuyoU+9EvodjaCw5ZTqZEsZ
9Q5eCsMTnWiuNV10YKbz9tvsVBgfuQ4u02Njbwhi8tuMdCEBCTJ7Ayw3dT1ANftwj3Sb4dma+LJK
o0ErUWMow/AF7kvfzR+TPUuGDCY9njJSt4qEAIHoz8Bf4zbRyIaO8MR0sUekwOxKS9t0kPPfzZ01
x2Ms+vI6Bi+8BIQ7EJ4vt/MhO9d4mYiPR1pmiqR8RrhpHQmqRpsStKfAPfvhv0wbxD/Qi1ko6DeN
u5sz28/KkgQsnKLz5p7eWuK7uOqep+iQQNysubLUgXs+GsQo1J2leg+3ayrvocWN/7APWCV8Gp3J
/dwavn42VBW/G9J+NOOB27nWg+TxUcM6N072Vo0TcxHFZ57eNUAiH2UE84kK74ionxsCYMgYujZu
5s1aTUzbLB3wdXdAkxEIVrFJ7htPwIGw6h8HBsg43YAs50SlbXbXfrYcindQaJYSuWIKk6iMkh5q
2qAnSZnHmPvBkECS8m1/0wEWXP1YodKfUp6TWxbIi2ZFI7PmZIoIqWdQw83eaiZpgrZL6Xr54XvK
b9dwuvy5XJLokJogjGyEefeb8plf1nUiiM+rWZm2zZ9kWUpPtbN5TgamJ/CFsI7ubYgmGrv+i4PF
rjOaLGZJ9CwfF8qeUX6LvvP6QCLnKv2tctH8PMB/OmkuuICFw/CCJ8rikRmIGuCYyi6SyCZWXmZF
bAu6aw85jjIGiGmYBvI96fS5o+0awDdZ60q/Bpc17xFrlBuXrdVmzy8GhWDsYH0/OCyXF4bCjSsQ
BxpRnNdMkIJvRMMdyrgYuVUuWmNEncxRX5A0ImcYylxMPXnctk7qorV+gNRImIIBnN1r16nSTRMs
yZIX1SfIn/J4KQX51u2N4cbigOOoIrKgso2d4ebFIHje4H5lI/YldGAB27wlItJ1f0Hw80LtzVpf
VmdG0ipvrC3i1vnqjNTT/UvnK+YIe9/eSoHAIZ5xrQ/RjptfN7QFEZSjJSe3eaXazidsR7YUs+4A
XE4Fvq+4C0/6WssCb1PaIHbbStLnJ/b3hl8G6ZTWObUwd/CiZaYsBYCldPF0Ki6YPId682TeL0En
13HZCOw/mz5LL9XsAePcn/QWJQdeS4K2/z2tJCAtpoxOijwwhOq6cClnV5SFN4isB361L8yE0vgg
bDHYuwWESTH2VTID+RByzPf50LlDgZXT9HR6rvB6NHAymnQKyKcpDgycXPy3izqAMuaDM+PN3UPc
sax5vPcwPg2epeD3L3VL/P/hr0Brp+P/Y7Kzw+ltz6R+sA+Z3Hj6upQz3lU3Qo/kKavHzTleFioA
xnJhAurIiiP3MmsLeVDMZJwmQ/osIXQ2IEn673hhmBK5IiNXqkpEBLZVFKM/npOvbX+Zs70+zkIU
1C/6BWVfJk4ZsLW0HHmV0rzIc13zOWWWrDlIQXDRk+3szSlO4SoiEHK908ZYqRc850qpFkf52MUn
nleKrhmVSHysTcZeB3iakRCTy4w1N4ZWLgf3iOO1OO71XbUimWBA6BtW/8EEv8Ju/zjPcLRF+q4h
p1yM3ypTNB6v6995PkxZdNj6tNE5ylCglLZaJtxqT09AsI8fqJ8lXtthUl89z8hfJl9f9KinF041
p2xjXL+2KnKrf5cDM0Xr4nyluou371GvUulWQLWGAR/0pV+sU2r4QMyb9qF6iwT+2yP1AFRfJGYd
raj8w5cZNOz4aO8JhDRKeeRG0XsiET6A1hVzNFFwL7WM+tdDSCZzThzsBK9Is39wN44ZXsg2oUmQ
yFzZDmEjnxLYmFEMJcngGW2qt+5aRbUcmKiuJD2skoC/USp4DKhm4t22syuXHaow3pf/6Xr4PG/b
auQe5GLdNIvoNjMYZ4Y0Pvz+SPAtU9W4ij6l6hsRY5vssDTzkqD91RJIXi5e9c5tMLDi8p2Am4qX
sXGzX4/BEMqLup3pS0uqzuK3amX2VELwNxiZgsiaiQCrg/J6L3qEavOIfGcW4H+jvHzSp0L3+/cc
7yEcajXdY15VmusX6nateK2pYEmADE4hGuA03jvblBGWrHZVARd3sT5laxY1NyRaQsRQWgc+FOJo
ALjBTAx2CiD4zehYpc4X1LFIQtg/dQXut5NZbBIDEqYD2TSgoFG0D0WsqnsgdUpvlKL7TGregvBw
G9PN6424Mw2uohDS54I5gZOjrUBAhSuACU4dZ9DD5jLFGXQb8Szyya2yU1vheSCbD6JY9yt3YBaj
M6ozbCsJ2PAOjTVkrYzK/nH65mIeeyVYZBr9hZhUvlDaJKQx/5UuAxPPJmVbgI+SuASzdy2Vhswk
L19xAOceBJYWnK619FumHmDAxCB9o7oEg32gD4kog+lsx0gAq2Lwn5vwl3IJm40UCnCd0nE+Z2rC
xwMThJyHK69M5MCakcivcClDx4PrfmjA4FSAa1qFXd1GPJabWz0QiF6VjflYW+i+1ONFFdFhVnw+
wVlb9rXbiOR50bdS5JBRpyycPWeUY06mhqht0cFqNd4kvInSe0fpfngzg0LurO3Ub65SlrkvIBQW
UARwmZJ/4zB2LO6VuKsf45w/wH38DS+2OcH+svDdwziycKsgNiUcV2s99DehPqpa07jgiURcAoZH
Cz5Cv0Ttnz7hKzXLhcutWSBBGG4Fo2oOhosHaOco5njr7LNzBnFoiTha32K2yGXtHpAEwrH5ako0
2YvWK4zUY8wb/9mm4W43jAqKOjl3NfXB/ZAivYMluM7EZJTYOPt7r01+Xo6fpRIjZLKB4VKOjxS5
KC84Hl+hxSJuRYts8UBAqyd1f1EgldZhjwrUGoarDHoDyFPXfj+ypuAJVd1HgesqYm2S2fzfx4bo
zh9WbhQkkL97p46pvmFb9wCa758OwHfwJT8laXC2lhuRG26lHYU8eZfZhAuj4ppoH3Gym+Y2nrz4
wZWRqcUMWPVz6OcDrST0Ka9qsAIuLlg+nDCBPTnXVVLce+bi1bIX0mFOwQuOTjS9jRix7N2CdlV9
KrCZv6Wn56Gi0ncv/wnes9W4hBgnqLE6Tk/2FsVM0sqTcq1ZFnmtX1b3mjS7In1MbEgHn3CL2PQT
qkeHQ0Mext5w7NuqvaBlKoHed0Thr3Bm9jyU/qm6cU/7ULYtemRYI4Si3KqsIume8tyBG3FnXVTB
moiYNpo8hzS8HISIil5KFMs+2WHk1jwXIlOQuX+MiLRoq8Dgp+9o+HC5j1hsg7JGW3araF149q8L
mBl/JQcOmJDMfxkjDVPwKK1YBT33ujbo69kAK9B5lnOAo1i07H8Rht15z2HEFguSmIb5E4/2mK7A
Z1WHwNTVdSkRbzlXIcsY4dzVAgLNFPub42JetSWjzMUKFWigCTEIdZddP9deSTTXxSG00ExrbwrO
lCS2v6oROdiPLG41NR5FwkW/eeS4F7tdP/Vjl1N7QLnu04JCfGrxuQI/o1ZHQhJ/dinGY5UVr+GA
YNLGLNM0zMmN0c7nQw6MGKCzcuJhFs8S5F1PiOIZm8/+Zx2WqBbISl4Cxigy0uk+EyVX4Jsdah44
SQw6MdAgZBow+D2j2DL6qTEOkv1UbIDP0pgNxoYPV6xSMaoPb17ESF8AO/omDQ1n6mJ3VveFL4zN
2NY491J8KQFTXsKR2+GOfJMT6Ilfe3HkVUHbAHBgcpisTXGWNuo13SPTxu1BhdNbqSJzSvhSnV8b
H3ng1+Mr71Jz2XDkyX1b7hHWyCBdY/oib1GQ8xFfUVr/LKJMkgHXg1kFVrHIkV+VvaMfMqw/Qwa9
v8L1XX56vS3ZNow0w/wKS3LYRlovL3HtKQXHY7wr1jzGLWuMlppYDx4I4jaOKtsrE8Tfxg9PUXje
AX/6B4GQBeIk1b0Yq6C4ffRynKIcSor67yOJWh8v7xupCSE1PYDNJb7HmE7zBC+T33w/E9vxQb/3
FIlpaskeIqbfVH7QDC2u13+GGvxT6J1oBcpkrGlWbk9jvt+VMhZbC3tewls9zlVlQy/TjBTRg6mn
Gkvzd9tMaM01rcPpJJbyMVYKWoZBN9d+13L0m42jqxSxEm4ME2igP+CHLSjHHHvEjUCxe4G16Zb3
060KAD0a0lqqOUEVu93bNynt1ehguU63owUKyGDt351+GbEiuKgQagTf/ptgUnsc+aq7z+nYty9p
VIOLdof8KnocWTIXymtjPhJ4IolTxUXhnoDZoD1/XY3ad5yf2zPbLgtFHeWcyBDYbYlB41RN/c1m
uMGlcKqF0ZjVqAk92G7TmR3jkn4eml7nipczz5KKwOZzFVAi8KdOxnL4btiBX+vx0JF8pdnXg2v5
a3XEQRM90MxM6AtaAbXfK1Kvbx96R2IjLvuXSAOlByplLUisqFJG6urxSDjABEMdg9wGRZqIGfVa
dGploCupDVCZruJ+0ex1gXoEjL4JH8cU1RVpd7MtN9IW9xZwkXv7Og4BPT20DFYgcdwC260XHSk6
Qpo9Ir3kH45pNQHQa28tPmMe+TLJqKjcLeo5v5s4grCVr2BrH6lhAqrWEU4V9lxmU9sAvP+0UKWw
9WzAEydELcRCMfqcFNad+YT/o0zxSI79x6G39HceahfmuFXUXf8QRVL7AkLo9MsYWbpBro0YUvxb
L9m4yVqA0v+8tVGGxOqNQ5e5iAJkfED3ZW8m3H0HlzfhMgR+LkFfKixpua1DtiwVEPuZ1Ww7bbGa
VkS2lZf0sSPwS/u3Yujl9OZ03ZPdEFNJKt7o3zwTG+JQVHc1b5OoqHXY0qPfK8POT6Y8P8YSTwwL
6ShJ1pprta6Fl5FXCBIptnj+MizyBXIcOmVPYXBlNnp7qkfFUjm343xJsMGDDTbfhLJCUGif1Clj
088yHATQfHiL45qKl7uS6WQgzobFLJo1IvWMXiXXMrkOcWQOQSia7uyZy8qtBCUi5tKU4pZRO62L
u7zDLPaPGfgu4BLPDYXbrCTFgbPX7PX7xRDIVN3LiIhOg2N/fv7mbumicdLchtKUTMecrzU8Orzl
+eXUqb4zRak+m8Pfmh0w9z55j7whVRGr7epMO0G6ARa66H5qio0UuYN/gJ+E5Kov8G+8+rJaEsqH
WasQ0+/ZZf8DOxu+bbful0/P70ZCvOehH3LymmKAYTnqg/JXYoQY7rqRA9CcwBnLB95INwYrhtGO
v+mkU+wXEIe+FSIlrE1adQglbr7A9IPocW9l9NgUp1x+t0c6wxM7qlTh2a1TqO7w9rQaJuDWhrgL
ophvt3gRoc5RlzSj4RGrwEKLHNf9AFZg1SagsWSqZ/DiOGOObaJ4G14WwoThmbJRwgdc85Z6dx9d
JbIHX/SsK9Jg65r0f0he3OwqMxI8ScBst4OXNDl4vPjhvUPbnFZPzKphhcLxNYC65AroKr/gDTRQ
5itxjmJ+qiUQEZLkUNhZH1qLBgOeUH15Cy+JsINkvo1Q3597DFz0gGhuFqVAGA3I1rcOXOjWCWb7
A3TxDxQr9UJKlgxQWl+7ye8C+vgaMDq3fzSpIRSbVb1YhEHBqsx5UGuJ0I1OpVKUw13L4DBso4Px
KQ6/HHTgiuK0UdlROEBPJBIUW4PmZxkqf0AysrD7MODcxwiNSqV99qWJLljvd96tJ/T+EbD8Rjxo
RHe9uksOAVJWgBxWmQXjjeEhvtgHcO+3c/uJmpmmjhuySvhK7Ji47j2KAWbD1mm9fo7fgHiVCQl7
n2slCPynWTcgK+W3JsLrGqYTj/fKUR2GGw1MDT7zWNX6/kA28yJfyIm6qjqEIxVqC7AzVw9HJWm5
8h+71bp+qPklX9mWDVAybZTXmjzQOmWV8NN9e2stWWQDE3XZ9pyoyE3P0Q8Bi3PeJ5mXtaAAzNdR
FDp1ZOk65B/apjXIQ+HMyjJkbiLtOtp/kXweHRoFIxCRElvHbkXHfjFNo8wbUwtSl8e6IaBYGUQr
XLIssw0aIEsd3wSyfOFvR6DvpY/DPmKo+ftWK2im8wUff9KBTmgpB8WgIcZFZxhlOLA9u+2/aTPT
PO0+n3HIw6Ei6NzWUYIXaQSefzxuLFe8uPw8awbD+eQH6MKqLdXBgsf2icZEE0Gl+MILPTjnCvl5
KKPltZrLCf+XhLQXCOpYsb+CD3WwuQCbsMQDo6NvsawKylecvqVTkmPgmRDDXkH6OiDZFfRqrDNK
pRMUqizp5zy5+nZV7NPiDxWb3l18Tariivn9mipgNBWZb2dDu5mbgYK8TY3DCzQT9qKV1MuM7x3W
9oaUDOpXnwsOImCTFgDybgLBcsMm/7Tmt/c1Uf1D3h/SzxTKKfKhGLvvZj8PVImej7Z24EaB6UFx
hPyZPCd4tFEI4m1Z6hE+nIFgWMVfGHTkGjcmqE4V9axfkOm2t+NCezfvsnwopbs+Z7GLDA8dFGar
5UUnjUIpkUqSYiQHbZQxqR1gGywXIyjsIJJTqcBZOaboy0GApbRgrdch2aDbYH4T3/RKZ/A6Kk3l
APDBQw0dIG+DSDkW+w6bs1MNhsXvHj0dBSeJAjbS9SczuetBbKIc9d/cAGGdu6OtuxPOGO06YZQK
b3ViAQSjvF2TFWd+nyUEhv0XKj85JJn+IlhpFvhAeI1eO5aI4OMBmt/0bIjKNxk1g0Wm6HSRoe6J
RYiCJT6hFGeyOGOyW1sWY2vUb9b+Zi4OHH4ipWkYsMw4rrubSZ/gbu+UnI9Ny1V2YciQNmx369Wo
fPtsWLUc5yVgVRSlmrOrDaNytMhnMNv7QmCYD6HKo6yPxsl3mba8UDWnueYUsOZwu4EmLd/p7plY
54Sm8xLLTHPipX6Vwv7UZ6SoxiFtVNMErlng+AHI8PNoiNI+pF92ALYnkFl+NiKlWZ3fqkPFGgC/
Fre7MQjK+iUhBfB6uJQexfWi54O4gDt+UImQhAJ+f4JsogAE+1vL+oSuawjMjrFAsQd88gEDE7x5
/cX4OeR1NBFLI80vHcWxDw22mLi3SkaSXLINVQMTNLIirJwp6I/H3YD1qYw/XzPa+AL/3OxNqh12
6KVdj9wuqO2uFZhjHT9xZCmff21szx7w7Q3TQj7oj/p9opbuqxgCKAbDDrCvdIrzPcCyKI0VKJEe
TAMc4uWTIwbC2p0y3zx388aTdzGT8+jFa5YvNd/s3oSRoq6Jg0fWQ2ydlV8sWcQ9u4CZRL7G3BaS
jhKUn26V/P9JbmyZCR/jW3Xf6zhmwHdfcFimiIiWqcINko+cKTS5G2PQTByl2t73+z/MwAjZ3QG3
IPuLu4aqwBXRvu8UQ40ldzpsRXBvLzKg5W7Ax0+2/TjOYoiaRlKyED5P2rKiIV8KoqdzT4s6LJ9x
2so8n3Bn7yBKvbvZv0kJUGZtfwqUDNhyBx2nzZkZX331Wzbj+/hrpzMnmyNQ1QCJq5ZXBP2L5ftF
OXZeZuUrqJFl6+eseeM11AOASXdJI7UW4zEswbpxmCXKzesju48iIjUqIrdDPSqbZxemkX/yqJnK
Xy7Vdo/DLcnJMTAOIA8wElNB3YkbK0RDJXH6ycAnqfsCb6s9k77KIu6O+ht1MUBn4Vqj0lhXWRGZ
MNraaN9IrCeyrZrQ6HTrqNn2lRsNeBvE9+00ymR1PzsugGHm9nnGl8Agw7O4ZqLIG2FBV5MSIKG1
9V8DumsKNAzejT7rT26dN38Wo1O7sNpVIXgiXg2kQeRmXa7J3lLIZPUNeGezxLhDJZBIAXn2j5Xj
cIYcWQ8VGD/81gtmTZnOVhmLL+r/D98JYwe+LrtzXujZAk+W9ViFtdt0W00se/DuNYEcpkXkRfMI
uDhUcDKdF3490btoIAng+HGH39FRi+DN8ZC5H6pfP2uTsvNoQaW5ol0+NW2oQzRA4zVeTel2l46Q
wSfR89YVMU7ow/wNELa7epJlSVCQA2il2lFEpvJ6G0LY+QgvK1z39PHFdqlivrTf+7dtnDYU4DOF
RLxlD51d5kpRk6arCKSWWTTWtBoHoKxdQaSdo2L9507p14sBUtzgF0uNGAinq96fvyK97BMYFUZg
jCr/Sg1isGIV4hUrr2NEIVZguCgEtW/5DDTVfrDfiKYCSCd9sOi6V9RFx9aNFuZ9lfKhGh3SyOYp
JxpyB7qP+x6o9F+Nabm+5Y4hrbUHofiecnJspf4fkfQJm04RIFGE7Glb1uUOBim8PBZaj4Lz8TDp
Qc0+7FYylOVeAPkBe4Xa13OlXddFJ/MeQOWExGoJha1AljuvYgC836orVRd4juMbmoEwAUVBRf8O
oxIbD7OaTabV/rHLljeKKNnNIKfPULLUmpfHUhOhbYGIpeqL3tYeW2akPQfr5SkcVnfQOGqfoZMi
s4Xz8zjPuhPXHJxtlPcsp8NQPKi2LYg6DjVBnsoyDZrWwEfc/gTu8Hyy8k2EcRsKW2T5Guyc8NI0
n0XCXvZNPmY1mkXFtKSvWzziFtYWkPlZZopQ2nFUFbcLY/AoGo5kXQ5VqxPZ+zH8+5vnSuriFwH6
HUUs4hxJ/m0VTtarZGa4qpvtzYjwFTkLYDBuSwT4V7zREydWEFjrqJRmJxljXKT8ljnfyFxJsgRJ
/9KbgIAXDKN3uaKrRIBdHFTzH+gb3XCiVj6BRbf7eNDKNbKW5v30Ui6qp6wJ/2OLuN6oqz7IpExg
ImFiCVEE9xmNrurMuf8byOdnCZUCw/R5fy7TX+3wrBDf7tau9PzkUkFa23O1pgrit+x8VbN/2kCy
PAi79DJvp5GF4pOdD8T1QYEQeXxmpI1zwrTcyZxoOPNsB7snJptq9kzkJnxO0PFJFywUDKAxprjB
hqmDMrJ3Hg9AaO+JkaLZKm21ZTSBEP31XeU2bjMME5wnfkJ10vCfS5ekqog8mBA2XVuTpqOAYAL+
Xe2I7sRqwUlm+vj16zuYa8nxgUg+/qB8cR+JrA71N46kItwi7jcrLOTcwSztR17FaYKa8ov+9eYt
W5CCz4L+DCruciD0YFpzF5vrhMDtXwqGJjyKD1EZtD5JUbKTKggjpQ2ESjSiMaJGF98+tFTDXsBw
wX6SqsrE9ZOJMqxmY9cZmoSaHySouQ3GVJ2IMwPVlxFRDSLiB4RJIKxbyukUi3FHqNfVSdOzAXYt
8ng0TiG2bw3K/aX7kqzZTvKMETsill/pjo6y2bdkN6Aa8082O7ZGAqA+MM3WRwUKbjboTQuHqwbw
0MrA1x8hgPRNScGL5h0539GuBXZ3bfZ5N1nDXFrMITKkM2aDIx/7mZC2s13I8pBPV2L4kNUtZaDf
wWM3O9jpT3RHOnJl0DTD+aESWC4CDHfnhRTtW5vy2F8ubnbVTPIsd1akX9LM0N9rMh9sdA/cUiw6
U2ZV2Om+jqsiBA9rzPWrJT8XfuubIp81uk1u8bVZO4fgKB5vl8R1uE5NHa9SqNJhAM03Tbq+qlyd
LgXqR2clcjTtFp662M0xX+zGkWndCVxzJrzXiF07iL9BRo2oA8TVl/eWORrYlq7/BF0N1Vu0rJfr
jb7AEDggIpuzXVAALWTWtrtpJyiyXt+NYIJM0qvOeHa4CoB2raH+3Pdhh0/XcULBMOjVWCWe1qUS
e6ZiHFMBsVPKYBYjJQUgISQ4CKHTkmLuWT9b4AqO1YqzaY7sSP0PFln9bbJeKtRGhCqwLk4h46gb
+wgk34lUFabku6McCxccgHdTfSWAPUhdVaTIZ8kzip2/+vp3LX+1ugwDJCtLTx46OhldiqzzvTzA
8PkwBCL8cfTjhEMSj5LWSm7n5NGRVy75DUO1IGAcU/cV441TIRTqYmxAOOF7/zLAWMlA+rfL8+kf
QbXsItW4m80n3QaKkDxS3pCKqghGWsHHBDQv+gHkTGiJjrvf7lXIYfzUiN9Ib6/99UqB5lZNhn3+
edctLfcKUyES0E19tAyH5xg9EQtRwXtdGhOLdS0ne23BMc+am56VoAffhrO4ISovZBBax6eKCZIA
78YcACr9ZHQ5bWcTm+qDyie/zYiInhz2nRg1o8iVmdLbhn+tL6JYhCr+A66Zu8tp/pZsCoHvtEMa
hNJX7ZvKG0gJNSgBlWb5vd9LM2qcY0Sb2LluVXFdGeCptxYYcMrzepFQGOmAsafp4RDKmyo/zzJV
RHGI6E6z7uzFgMUR1P3xPGB2rN+N7Wddqlcn4gMWYBmdRbalUI6ZnB3HYS+4y91QwFJKR50nv/R6
oZrfToTA62eFjVuDC8z8moCGR0rE/38nNDSIwqORVfqAgW/GUJIZY1YYeHUksMoYuy/uOaFfmmSY
6C4LbmTr1FeOpadAIetz8JIOa18DK6TwQUQY9LVqeZ5uMOogsmUOWWAbNRG0ss4ABk6LWRTD3soL
Oh3BURRN8DnU/UVsS8daPax3UxvJernczQDN54TvylTArVaAsjrdANjoq9LP6Y/CC41Otb8koNML
dCudrZBnP3TzXsxqE8hOlBk/8WUXY1dZ+scVKYV2BcYUqFojKn054Kb2ZszyrKbrU0ynDxWEAmhD
rzUbJsZNaEAQsE8bStOSCAyC4vzut6dztqbLlslw41u3zCuuiUdsNuk6DNg2DRr58v/6NTj13tBH
8RKnpnI3jfccOGeBz1IHwiWXT4VgT90PTXdKseqHX/7ble/DiPuDpAJMSGUvJe3xfgsyMr3rzNek
WjZFb/cu89ySKlamjUGIKPw4M8otsvLDzBX+AhNC0d7mKZ6w0HweOlHDPln2lg5uY31Zz+tgMIcw
CgpdEi4EdElp86SDUaLBZ6GcPsVXuDncoVF1JqY8ehKA6D+hQBwBPANNOZ5pCRoCNR3kWDV/jkSo
kVfvrKmG92etEkP+SUOausad7kEJB7UVTLHzydUQwzxm8pEql9nyuRkoJ+yoDid9Il9gQku4Y3W8
v06vonpOrws24Z7imvx8jerxX/I4Ox1FrAU75kbVLwTN6bmGax5IArz2ilG2B9ic0FbblzIL5QVT
jCFouYmEyo5BhdLYBkqSsyfW05K8gY/MxM5NJFX0qKcB2QwjcjtYTcR6il3SnxL0GUloNYeVxtxB
8ZEgFQ5dm27PgGt0h5HBCQF8pArQrTSpJ+zPpi5vEY9ZPledoY7ar996Sk5WrGXuBI9pt5kPOFUq
vAd1gT25ngxC7XM73B9SfTXkDtrTOGUoBY2wslIKsLUeMK12Ru4lb0J78hPZzEdtHNaZPwaGgIsR
AiDiQ/azWHKSgKccgqBg6+Ibep0qHO6CF3aAgJcCpwpKmHIzB9/rHoN4znrE4LFZecu2qjdu223P
TTsYZhSTkS7hO6ROSMc3HVphw5tWNmEdQAYfJMLbx7Ki9C9FNGs2gFsf8MysHki4E22LAz5HSgDr
56kiAy4isWPE8bkiLkw/Llmh9TjXG2MZQ5GdAMhIaTIpDxJ/+9NjDaWh7Y677dQgsf1b1osr6cbi
7v+HvLapklZUfnvvdcRqfPWNVINd+p58oVDpg5Jmkwspde9LjKwh4KOgMd2UTAiae0CKIpD8FewD
TaX834Ax/bQMrKJRaU9S2G80v/at8KyrsArbF6eUr8PzjEW5vL8Qquy9aDYQmXTlOa9DBwwYc0m8
p3pKYTla5TCPJlN8I9LKGNiGDvP6hBe1tNpygrvZUi7LFEXc8hlyrkLjbQUBHds/wseWqOTWmlMy
lUjI24l5tsLI4dx6ZQP+OmJdZ7B4OLui6108ZQPfBmqZQGfSBvE7AEjiiKbyB73sBphUIRqvsWw0
gR9xQk7Wrx/Aaa5PLqDwxszuSbZ5jHmkuwCBCdlWQGm6fP+KaFFKh4/vykCNn9YPxEBcOIkvSBfQ
+mlRovCGogzlS26sFa6uJPzxudng0EJARyUzkQQHFU/T5OIZvLq9Rv7kZkf9BoBZvUhw0O1jCkzm
zs/CmPaseLEokRoWthePeP2JEOLSUJWWgvqDwm7YZTj85U6/r32+ROtzU6ZjSNAcS8XjzbCKIbL9
YPUWkyYHjaVulHc/NpuiOy01EKPqlk4snENALIkDKntWC7nMSbS69lowoqBHpRlgYWjR5K3hsvj2
t++x5dRG55L/GDDt+dhNtWBoaaoaXCk3nzXcB9NsUYAA1L4cCopjEa086KaByNRxB9ZFSfje1CZU
ZSaAzQUe/ey57DSlqQTXEOjeUDVda5Vfpb0ZFqNs0bJphiXZt8smQXdiJbJsjdqzMwBfdzThAGZ5
OAO1+pf1GzZGiT7a5z6WEDFIS8u5m5I8AyooXrDGSFFjxJizU15Pck5Mpx93C07+Db6CzuX3VYS/
HHgRKX0Lbt5diruPzLsNQ0RNKtH11XUX8qLMmcvZC6yr9inGnkdtLJ83k/2SHIXl9nOTTR7PdfF2
DBnuBXM8OGlbrhzHkWOxUZlsL6u5QEGLW1H8rhpbG7V7og7TFCFPFGZbyYigQlamLUJJ+hkdE26a
AB/zYZSFd8KP3CGXwoTWPSHsgls8Q+rWneVgiVPGXnlO8lenLMqOzef+31iL21SJNGpvDX9CZo/m
eUB6TCR4L1KgOGo+ivkE1Y8owgfe1mq7P1FUgwuQnIepiuqIJtrGDK3giDn+cHr5nOMlc2k6EtG+
Hyncv17D03gJGeHa8o6JfG7z5P85eXL814iWAEieMTHbskJvIHw7fOBn7sYIXq9y9dfv5x1lVdhf
GUS53F6Es28932Mtet3ZWaz1McaYQMeiyXfIam0obVOFigGfTTjrNauJfWK+/RYG1wZ7wNO2NC4A
i7/R2RIQ/EzIyl9KmYrPDbZAHb4fzYHnMAGaj20U17j2ne8oX/mpPMM6esOF6UgyBp0SGBcOGjP4
HFjeLWZGwLQ0+0eJa7XSlBs87pqVjAxQboey0zq/s3GlotjuR55fWEaja3gih9lQbwCmEyux1qgd
LZVixUV/iaM6M63aCG7bcV7zHpIkamx3/xSNKjb/fIujPR4Elo6EmK5zxs72SvrY1NJUB3Kk/SgI
wG4oSgvGGuT4otaLhM8wCttS6CBg0QQYYcxyMqfb5aaF/Z978x181bv32+hzpoEXQYyy9+w2pVY8
cpGZKF6xJJuEOD7fLYzDLOO8PJYoiYXC8/LZ6rT5VQUFctpV341zdqqA+XXh4n850Ly7BJvsQkFm
7+YVTegMZsGunYNgFIlloJhVuLgpjj4v2oY7YFNQJORuLsg0Cv3rzG2tNq2CQRJBDKXcRse6TiW8
fExRfYdWwOYLCcXMTrM1Wf5m9bXEgusKAGPAM2d6uGEG55T3Dnxcdyqs9wg53CwzHRPelhWsXA5r
RFy4d4gZu00dmv82JXcOKScud6APJOVwz/Evh9Ua51mDMz7zbISF0TjK1pyDieLJCYdRsFmubYFV
5FwqpUdiKo60KwYMcAnMjg18oVPwf68flpdJe/KE4vXOJYpnfOH5vZhVjATNulEd0IOxbJl9jCWK
kM7XDv3nyvDbIB6n3djmHs0zMuLYeiN+aPb3Lcqp2L3NlpKBq/gM7wBDNYhG9serzllMjA25t746
eoW3idbiMA1puqM1M0w+fZ7hdZ4x6MHoRHs8hnvT119cN06IcOmpdQDwxMTw0XSGqUA8TyX2zxkA
fp+GK22uUwKR4eF+L+uouuFNYNPagZZt2pp3FyKAvjovHOnV0mfb229A6UrDUjP/LLlAUL5zZPgE
m/sVtsWUuL+fJX00ueNAjnZahD55LMFxG8KLoOE8fAmPEUKLxD92l1No//wG5LojQwu+YNL7lsp/
sufQVUi9mH97QgUPPrx0VbkxQxnWxErFLFNC9ammRGsrsJbUqzwAS7+GKpsAak0J+6P9j5AD6Iti
hWeO8GmdzcFR3HTedjQ2mQx1mxg7Gb2tgNLCBMw1Gxpzeu47yWELAw3YEPuIRqejZZm/bGt5cC8+
cDIrUzsrkVzSOwSIZuyd5uDtccXNuw5R2vnvGw+OYlDS93FuYX33R5sHPlS/uQ0vcpd3lNVcNBU2
SCyGqz8sHchSaKLcqrq2KjrGseZvleXM2sXQG6nNQp4VG8JIdFwreT3l6rBpWj2l7PO/FPp5KjTl
qruIPMaPDf72ebRe59ALbUpJ8v2A7rnzPVd3HMxpI526tXrD81Szi6TZfKbX+y56+/NQUYExEPtj
R3ge+y7Vc/dCNiyLwBcaTG2fqeRty/4ypTPCmx4rMcPAcq4bsOwPVHhEKJFRiO00CbOFpcD7WuJ8
Ohpgandblp8K/I6tTnrwPTZY0KaFtJ48mP0Zb9km2kTNftrnm/6QB1VNfF0jd65FfWY4rjLFuPbJ
6v61XyKTcTsu7SSxZlFH3Hh4DKiY5WaguFDc0laevdpWiePjqxDo4eAI7xtjtZDo79GNVjO5Z6bG
KS/uADtKdGcj8xgQrAX1QkIl8rtu3nEQN5mhZqyL0eseClbTcObTfDwdI+BbxjLQ0oh9W9O+UdTd
pVXkMXZfWLXRrzGwg9Tw/M5K+4n7oPVmzzM6UAH4CwbJlSXfDz5nqT4zcNsJxnOAN6HfMpJ4oLjQ
9m83OAq3tA/WzQYdtpSMZZZ+eyei0XTLDmo8NYttFEJIe5UK+JaqGBAtWj3rNlo0yf4vdHdoQnXL
Lp1VfHQ9ybe1KwaIzAfp4ChnuXPuJ+uXcmwnS+u558IZe+9l6J/UViXRstL79I1z4MkxRC9ypdd8
jbnBUc20hHN9nHjzB/x5D7vLug4SGtuyN8tsGX0Ag9qgbxo1/fstFEGtyFR7jukgQNFSZqQMW95j
djd2y0X2QQSlhU77tVFrvMPScN7jAWNGsf9HrLEytBsMYcRSDO1BGfbJyoJkYlm6Mkcd0w0hDdzE
ZTUtGnR83eogv8AWKsNmFyK6J9AnQxnA/VNVm7qpuUVxrsKH16kk//kxB25Boen7rzR4iA3LSiC2
xThSuVPSZtRgQGQdGWHmX8cnMJLG8bKdYkvEnYLwGet1pclbUZjK3IMZ3KsmL2nVK68mfRsxq51T
+FO/Owc3IuUrcwBiVKZtzj5vGCyPsZzFV0wn+wWvpU9o/aKwQahAXFegx3yhXznSqWyStud9m2th
QIKFLen9/k+KN3pwob9vYcTmcGhK3BGKKwALFnplteREPw7+OQOGtqb1ltZxgYHWGiuCvMxQSz8q
H0Mttwom8+IpKmQK5tbxlzBqJgVlfoU2HHfoJ2RBOXL+U+BZBsHZqQUgJCJI6QW+brLUkjUvG8Jo
26vV6F79o9oS2ld99EJHNY/y2r68h2W6YK+F5r00H5bIBHDPzHAmLAGeYBKnZVPg33mZ8nVCCzIb
5ct7PBc4var8QIGIBoMgn4KyIS4iLG9Bwl/1ypbKHRJIi/FwiRii0dMG4bBPHVAPKffud3eJsrm6
igAJ8vyYOMZqzl8YcqIKgqTDT0/7ZLoENnZLezrtVau52XLHgVdcxG84uFeANMjiz/EWH1XW78KY
+VW1vsDdOp+BnDBdd08xnnMBQ+uMNxuZNO7z34tjglA3pWr/e0ogi4JuKtpuF6BOUhM94a2PTvOj
2kzcPqBFZkKDsWIhGC5NvF3yRdujlkjVtLfDKbT5x4IJzRBN2yuRNYlQBjstOrr+AB+KMG5Z8bzG
pKBMOEwLLNxbLKJXFU24J+UkGE8/Aau7aLZ5Soq5JqEr7fgHjOSODvzdqwbTpH7Pn9Gg6FNc9sRF
1gSZe8Wd9T4wYKK2i1DbJJgXT9SCks+aFqTGpHfOE280CrgxvDvlgyKPs8j32rORtzn7Xina9sM7
xgnaCTdKQY1f4ky+zTNlaMVWSjnCTthkeBlkGrlX3MFBIATJd5fE2teO3lskUt5SX0fVxC0DJ3rO
Y3WDqDXcTNdUdME0jmVqPuXcDaOOC1jlRS8fn4OY2We66c4O93sY6KvKiSGqxcv1WRUAFuQWoEbo
wtOI/6FCN17peeJd8EUy4RxSJiVOWQ7sWh6dWAF8IoXsM8nqheMwf0WFAacam/UW0gT3tTG7yXvs
Nw3wOyN9Qdjyzz2ODRRAEFH/1T+1fI8hkg1bbmtsCfIJQDMUyOdD7oGRkWvkVkHjyfZfeL5hiIEg
1nrLNGe9hWBGpxB0WiGMbeu2o0AcfdDjjgo7El9lIxR+jOZ9pcfgXutJ83guvQYfe9lT2n95bojt
3+zL0abpIhvyil/SqSLr5r9K0g5jcMiUMK7iF10vBD4dVPS1sFEeZMUamC7Z5chxwdkE3lFggTWI
uPMQRXgUZ/XidabCO5q75r79u6rc1aCQSl/qAvMq3kM5JR6t0nyB+p6K1xocxlVGu7hn+saBTYCR
EUulqtHFkNXIGJ1GKXqCqxTedgdmagHdiRLZdie80Ij0l6xih3bRbLXHmIRmnU0c8uBrnOgoi8iU
ZtPeo9Z9O8TtqaqQF7Cjn/CQpumg5QZ/eL4nVUhN37gtgWkTUYwG9gDnZXadMBmW0E05FJRbrpd8
OgAGlljSoyYqgPjB3gOp92/N5TTwBO9UWKkWTjH0Xb+8Zijp+tgPz4CjSuPPRky9TpKC8z7Obwyp
M81UVMYN8+4KaBu9rgZpHVtDXQStpNQZel/kuyi3WZ15b/fmFsr4p+AxERkCrzt8gi7TOgcyVxSn
O2UdMCB2nj+ZE1VCriyRIfu2r4fYJPp+yS0tcL/vRN+y+E/t1LJcBu5Q8O7K+kZABvpDDvxP7AwZ
6WjgRnmEpvtgwoC3qSF2GAg6iaEpfmDKZgDkMvXTSz4zaS5wzC2CxI3BAlMvxjHVNoNBLe+hJaA8
mBjauiF/ejTPoTJiP+D1nv6yxM+8tIpsnVSX41IC2/FUxJuOvozu1GRVoMK41BIExwCbga2spgZE
Y+eju3IwqvgneuwSRyaufN9nXYPl01jPDwFlPSeG8uosqOr9KpghWXOOqOi531Oz8hGBUPLGpzFo
HU4xynUxL6kw8X+gr+S9yBqYipUU27ua7SNxLGxAaxrkX2H2//IQFJ7rjh0Y8iFSzV4iIAWh6mZI
0UH4ETbFKEgYhCUgS2l/0KpNU9I696aamHt8YhpyVyNS40HuZCdh9BfU0B7wcKZn9T4KcxhKGy5y
UFOJDZP/AXtxbue9hqycev/IxR7+9Zo3Fjchf5BGBo7nLPFMeNBEO+dxcleSoeAMZLGqIbIfnEFT
iOPzHxWCAgfN61WM2io86FDqTqgxxFE19TGWGhDsFIwMFJVrTB2yqwhCkQmJQUm7d7OaxOyFDGd8
usPVCQs9d3E33dMA81HfUWCls8udK+37CXJFd1z2uOzUDIU4DepL9S9EFgvbQTwR926hUVmHD51w
4rdW2Wgh7rT5SzSTkCmSivKv3NCn+XQeis8iEGhx7kDFNTOQZ02sdGd9RkZF3cbMQcomX+d+O2eZ
RtSLfyA9ofZ2L7nToABmrpO1dmIX3ayGkMMIPpii0eE8fbiwzcrNLn0/QfySJ0nu+Svlq/K57mWI
i79kvA0NP7+X/Rof+E2XwVFCjxPaRtgVb1qG4d+s4gXyLfxzRlY6/EA1X/z8l0gO6UeEpbxFpcCW
/ppD3mXPRW7v49nUmZ+kA+bqVbGTW+pJK71rcMpqQi2ZTr5WY3I/6Vw883uUmqbcs2DHQOWuTdxz
dA2HgHmxC1x6ds6aWEYJ4VWNG/eEbt2Xp9uHbfnWkUOcpRe4pRmAg7d0ykZvp/QKqUbU/y3vSzHR
WxhPDjL6DXY8riIWn/tWenX9DK18sJaBOA/IhTGm0CWT1iPwrcVNgiowPY3FQJ3y7xo8hug0qs8j
1e59VeqiSSmlOw5gxSxhaCzvV1a2hlLmDIKukzdVhILSoM805mdveY7lzJs5DbYFJATFC7vUpbeV
s4PwJFZM/M1hsUwiXG44suL2KP5QHr/ELerSR+MyOUn3h/PACnW7BQT1BR7RJzHD4GYewgY36QSR
f7qdrc/Xqk3oJ68Aw6SQoDGp2Kj3KamwKCw8rXpqFZ7Q/fcHRTzSGWs80+cs5QBLLuAbdNKBR9lP
+3Z4vA9nWf+2OOja7Szgy7F9hAsDcFZJ9Li0sJU9EbpTHg/gYtQGbMPu9mJbXAUj42mDMbUGEYif
aTKLLE3nBJE+OaGe4zyAU1Ze+zDe7K7Lh+VlfYzOvsec/BKGHfLKy0W86nyU9gqIIo3FTeVbGWsg
CmdJRP77A4q3EfCszr6aW1ekZtjqhgOwfZdo7naik1b1oMzrslIbemJZWaShIzPn9zZhqKmuBnEe
DmHNAPXzUr7x9NoQI0rSuLgp+ksth5b7XV4iwU4bqPP9EWvcFE7/KASgPWKl1GYyu2yzCNsr1xZn
c/uJWe2Dv/26RFz6RfzocZrrB0lUv92NmXDrBT+pMfTqPOF+jxyNnpdUojBRDjVPTaMaZtG83xLo
QO8tOMjlK/8xXhTlVBacSTKGw2wZ0o7VxNRd5db2FEe9wjk1+GKNgc45k9uh7NEJ2snbFu4fPbJz
6jEfjEarAmSjpcoq3gSFOLMAKmiC2cXXJW44c3zQQQbGoGAapTctu6W3Xy3+ugKOWbBehpBSUw1U
VuuzMzVVupYCDRXkln07BbhtkJkVREYB6ID+RlH2j+3KPpW9JKBxlW6qB7h18ONisk60EmUKSsTT
lHTgqVmQSHqPAcJo9yCVRtsrQkDt1z03JB+hN4i+ZFljmK8ENGtJq1c/lYvvyzQBg/nJQkQwm+P2
rDaXP3IDjFyL6uXGnIkqGNuy8mjQzjEYoWvpVg79c4/LRMl0LwfN5LAN/67AeaEDmzyyafe/iEJC
n5BQKFndptLTTiuCfCEdNPOQiOQIhLM9xIJK/gQJxfh/8c98HHLByPAXuHQ/xUBICunVI0YDNjaA
gyls4q662wPvS4txgSK4aAqpOH4zMVfW3mUKfZX+iKNxVfgj2qW3ATzmwcinrfwNY+w3sQOVHYXC
aDjqvoyLGOClYIhRRFF9KJ0qYx5vU8hv0kM/W0zUV0ZQ5IE42+HhbYbLw3znkbupVENchxvDS3Hx
NRXF55wJx9HZ4QSkWKUyqNgLlFGMdjGxghKf2vI5n2Bb4V7a0JpzaYmqBlW66Wh0cNl64JjVKG3e
jYDm6K+gJzqkgfdP9RveCDB5oDHFOIwdEuHaP4noqMvHMvEIwjEOls2j6M5lue3myPCRd6RuDPgb
7rmdzLAk9iQntRTqs8mcWm+M5k3iiqyCvnVqmbZzTe9UFcfwKsp47aloXFbTHtvTWBhvMqMQbPji
I0O3ZyWpzgFiTjwFfULDF1Abt9KKY3CK/xUqNWeYdNnAG37yvfehQgg393iGInArILJgzEfp7m0x
dZ7bOnAoaMYGa4xoPptTN0Zlw8skH9WjwGjyMvWJjOCuQp0OW44uYLAXxAk+inqiCgUzp0zddiuZ
KH2O5GBQdakWVx0wb8SGIexwTPAZee8zNB4rVsT9IvfE6cf8U3//NgSp4VE3V7OotNqL5elPfS/+
RwQ7Un6Pv5inO9gTYHz/vJrOfN+8fmOy+iPvItZmgBUcCut6ejn7a96hf93K795AsytfEi/9GM1i
SLlYvc8fsMV9+4CTQGIXISUxbhByMO0g892lMtCnY1UDaEvSYZ7tg+u4ZTHY76Ykg0nfOBq4UOVp
ByMdZTEemEF32iltNJ+Q5eRh4Tz9Um0i6geJBgxjloC4aEuid9wLLT6+jiEeKJaK5v1bKnrEIACM
yZNSLSm3vw491mr3jdScoC1cVQB4sK1Kq2cRvmoQTgoj8VwxlgT+DlNyTQF4Ya5x6/BLJz9WswRl
AqfTWdH99FV+skJFcylN+SAjwNp2dW2c+vAP7cOeUwXLWq4IWrvJY6qTi85v2MC+P2PRGDbIfLhn
Z32erMp2QTMuO2fLDxvjuSZBJ0uAAQSBJarako+gawstyDbe9883tofBDiSjqIuPXBpTmu/cyil7
X4biABCskWGHa8bT49mR2PEYYCQZ/58VXp3a2stw86KZbimoFLOndqvMTs4B8/v4Skg3HAxStdI5
Rn45BrJXhJboNxdgKjECWAGX3oo1EGLQI+/brMBqvg9UBPNUl9aMsn/wvclGnJlbmBj54cEHFQK3
FFgn4A2807wl8WulhyuLM/in8B+xJUoS4N7QjPaPr+BG+kazf/aOJ5kRTqvChd9XlFXCVZpZrpRF
L8/hmEpTsPuI/9wGUapUtjphJTdYjPte+20qj2pfGdQpvRJR3kcrN57E7oMvyyJy7uodwKcu1ssC
mS1SC8f+gBSN4lGtTaKNfRaDuDRq8kwAPoPnJVTXiRXLdXig0JfviXmVogd8/T8ia8lHqQKsv7qQ
6gFfVbhNnLXAN6OXx5yJtDV8PSFHWN7+DZ0fqtS/kd1PgqmyZiW7m5NA6CxHZwx/q68Fc6oF999y
ZhS2WRScRNN52bMCwYAj8QcF3uP4PCfMeT2lyJJKX45KEXuPHsNAEAkr6J0XLGohyd1SapuC5IV+
5CgSfgaERvnJt1ndX9rYag+lnL9f/2oQZCsChcYlIYRtp2FL+wMmw11zSDwPLi+rxdoI94/3j797
fDGfODVFxXw5+V2XIgVlTFttICyQYyX07I4mEzlnSyEQv/kSaX4RoaQzNwTBoc4sLZT90VIXUPtU
m9YVjbBWezpAeaXBc1xJ0ecDgbQ8UxU9OLVLI/Afd0GxPcpwiPvMKjfRxqNoFGwqVKubjgbbnT8a
6WE+w18T10JF8LiVAVsh/Rq72QXHdRyYrbPeEZACajl5WPbzDcpxor5grYiIAu1uisZyBhQ7kk74
diizKGxkaZVavnkjmPdGbZrr8ESnB/1zG9JmJRxbo5anT85JycPIBWTmepsBOsQn03YKm339Ytcp
88yZrK/+cn9N9niyO6en6aA+tkPppoXUpY6TD6A0xC5bEH5oMEq/CvZYmBvBeeUmMbQ8OxekXjcD
hTAt8fdvV23kxUtctwkBfKiJ0AXmzecTT/3IGCSgvsvYJlcDqQT7yub3Pc8ncEW6EOE1lImFALO0
bfxO3PIDt5ZnXGfN9qI/C/xtsd2En9aXngY2qOFw/P3dZpRJVPPXHOUe2seEB4jq3QJhiPcsF/x9
y1iImPK+EizkJLiZd0ecrQnI4BALoazNg9yXndcgkkZSo+MCGaN74Xvk7YdMVzpNw5cG8RdwmKXA
VaDz8g2FhiHfjPGMKPAsEYiIA5Eblih1XDVTp2t5vUzbk1S5z9XUvySKTDAlkAqWIbt7qBsdnXCj
46X3nSB9IQtl4h4Cv9J1Va/E+6f1RcKnYejegR971THVSD5/RhPZ5jrf7FKHdzGb1M4LOpX3Dx5x
3rnaOwFR4gh6mxH2mTHaHvYL9fhNGG6H8rYgZjcknsUz6UQN1h7w5LEZyEWI+n693esJbuq6v/sS
kO3fjwZBMdgaSb4g+bTceU3UZVGHlrB/2c/i9uxvIVkfSpwWMUl0O7kYmTq3U36htBuLBrm1UFnC
9d9zGz/82s+XmJ/bCiTFJqyH1HUfHyhx9xIcXQrHDjCytaW3hOWg7V2F9DvU987AWO/bC26Fx0Xp
DxgJ48+6Z95hg/QhhURckFKd1sJMNY9zAK8bdn5K0FgTDfjoKiMi4DMUxlm29F8tkjvvcGnaNLsN
n3ntmBVMFlAestFff0FuzIU7XscPqGbp2tZB2Z8tESnXcUCdmCV35xA82Z+FwNpsln9J0qjGoyZb
1FOwA6oF0xMV9harDt8FKckgEkV1XkYVGaQJwGdntY5ajQwcE13Szh3lP5mlW2+OBsU6MEtzWIao
6CoM7wEq79jWISc3CXQ1at13XD7XvTseNNg1lQa3xG4Q0TENfvjIVqwVvWKrjlh8jh13myje2P93
5QGm0ZpA2SqFqs8WJOjZQ+ed+H3qt0zS13CSNuvmHyc3g+BH7GIJb2rJxvCOhQLRHIvlkTlO1Ac2
W0eoVM9KhxQBnSJlvV78DcgJFBUQ+OJR2tlvC99sZ9oMzAQNr83NKOpEzXDNyTJA5j8uVIKsYRF3
w24k+aqeIlIbTK/ahKiE9HmxMHY9sfyGUdGEU1nawqoZRA9WKuHOmzlZRL+eHPqlyjenRuvGTIXF
Y7G3kf2gY5nugAZ6kngj6Vd+ekqLd3YkOc//D+6iOERc2Me+o+ZK7EZwtZ+UkjxVlxJI11UTLswP
guxVLrTtvwt1RUpUSKR7mevac182B4MtaxEnwhxx9BK9hlaOZQBvlLQchydm3Ttjye1KC3oXzczH
zU/ItfVpbfAN7WYQNBTXunUmNeZAH7AOHiLC93vOhxnrnH/AHr2F9xB4IMSpQPsdTjI0gjWPD3QG
CUFs7KD0ATy9D6JCcr0kMIy0lIdgjN/8jQ6rMPheL8Bw7wVWUDwbLwFFkzX1oACOdQkSenBv3lcS
QPowCqEr/4FzrGl3iYxXsPQ40fRSzBTid9I+12lNI76MIZ8jGNr0rRWVp/6echunNGmSHGyyP2AB
9h5qFKSW479++tcLQtyqDSRMG2udfQtTzCn60WLk0MhIRg82RHxS8HxjL5bZZvVAx3PiAWzh7/pV
QeTCUyep/PlYgb6qQOOlwLAtRtM7n6GZkEpXSyHXInYfTnE3wSoIgPLxcq+9NKF2gJQDeBXv+gEU
rIdGavPBHTX+tazPzqgKl46x9yMK1UT1vMY+ilVs5VfShPYx7x/alWP+x6+7+qnPA80outVaTrU8
1C4QmTg/gIHbxXPbdljcUyZBGIN4SLRrjVOaQ4Jko479aFKTtcJG8GbSWskNw7m2OpgGW2smMH5M
0G7qto1jidiH26wtD8qpjXTxaznjYJS6GhKHrL+jymMty8nNURj8PuMmcoI7Gqte3zhq10WzpxWW
OGhSjU94j+jzdrhvNYLeofu0wb3ogi7FWiU6x/fyiuar2gNV5q5760fX+yE0GyzbWW1MuEeArKvI
weTz8IAEZJYzaojVEnfKa82xBizCJjg3AHm/Xch1u/ML7x0koESQGS1qtzc4O4W5WRRfw4nukd69
xdvtTaDHllU3pA2fmGj4Bgq9B9ybvW0XJ64iJc87L2chvuBC5dHzsJRyeXG9VZRqO/CpxxaFeigv
vWdt8OCHzUjHVHbVXrif4ZpPJTQaetJRgX0oFNE6IFsNOkL/aDF8vS4CwMpz0w6r00AxUeqMvDgi
vKcZUrwf5rAp8j6u+CoyoYyflmse631SfGkoZhehayRjcbE0EeLBvjsPMMNx/k02oLaivLxR1iob
/3BYsEWadbAW38sDMDuK2X+26nGe7VWYfLyngpdh8scSrKDQQlxixP1byzoOSRqhwKIxPlRBW1fK
wpDSHLQXUdd/90I12Q5vnHL8RuleBGvkiyqmleV2Tw+lHXopB2TuTsqH4hXLQy3B+z3MUbd+GZRU
Cnv3uu+aIQ+2e43zOPRBpKlUHNvydsSo1vCMi1TA8F3LPs75Op+aB3wuDahdQ8dfKQLDA4KmO+y1
kwlDMyLecnSLw8HR+MVKcgVx6BaRpqP38gX5w/AW9aWJZVu2y2PsgYJ7o+HAulnT29cyCCNODXlJ
T763WLSz+8SqJ0ZNgpd2BiP8Gp1VqOzReoVhvD/XRDBq06RHoekA93F0/HCe7iZREWVbtJy/sYDl
/cdg/+iWpHmuxWfR2SuMiFc8MZAW4LnOo4i/7s4WVEu9Hg/HHeP/43gvh6l9XfrV0KhYIYBuPZjw
0RClTzqfpdDGfvisy3SI73fwaid7CDgkoietI/O3ozl4NWU6k7oiH2tdjOfwRzBtQxouaMtDN0ZP
A/qPWj2l3Be/0IyrRzMe/M66Pd1+1RRrAe/XFvJuY283TgFfFiUds7zX/a4AOl935ePiPUklRe8t
QvhpiqnLcIeCQVWDPQsg0q9lzZlAqhm/7W6UcpO5ft3IEcgUnpnNXbJICjxS0c3RRtxZhqVaMnuy
2PtCBYXL6flK2U5Qfh4SUA6r+C/kF8y+VPGJp7qd1A/tgvsJXOC1or4BZP32objRSg5tI7T90dCP
qyc0iLmuYrOD0rO5Xxape2y/bLQTBZwJZeT+3WIWLHtwpy6gKoLjol3qhxNdOYGPn0t9wI99CH1+
V7CXiWaTiiaRZV0knf6F9x7qEkUS5T8njNajg0yVecPmACKtorVh9BceGwsccj+mciIBymMcTZyp
eTPNb/6o1dG8h1ZkZ4ihhqILuY10hDvHW7mqS5GKi6QHxhnSdT69Ejy1pUQUoUoXr/Y7UeYCP4XL
5NdtM1F2FaCsEWilKUcONEq4LvB4jjh/mrmNJKKqVvnIN/AJk57yQO9dpSU4eYvG4mE+SHCg6eUP
c6eaQkvcJr2ycX2ivB1UzqxfUMtRkgAbt9dl3efybi7Yj4LppSzBUYiQ1SHPJogBS8Y94jlAlGXt
8GEmI5Y5ydO1fa6hM0sNS8lERyHO0moqGU2P++w8h+KFv00NbYofqEkmANMuIul32wyTxymzGJ5e
e8Kyk6Uc8s2RqrBCDsaw5er0+jmwkKFB3DNMfYgnp/lySuDKr9ltNHw4gkgycNhpT5FnGqlegqCs
qyWrvupLQVZ0jB1uZwg9yl0QCQ3tRhrmr6ufdCm9MZDKJy3+QGr5Q66SLCCV1ycJERMn5mfBnRZj
nJoM4ETzpekJKMUMurvmEezXAltIuY9x52Sq8LBMhSIcAMkJwp0a37fL8zUFz7Lp2YjuhimjSG0O
izCsnCWLs0ZhyX9qw+CkSkHGf5UhTjRTLd5WE6Q8AwirR7MefDxtKy+GkVe7JNcMN07HcfNERsZo
uh6NyENLDtSV16VRlChKeF9+FQeZnSgG/dnggOLlLhr4IRyBqJt4vMX7zd2vy7RDNtTPZ9dsQf8L
YiDxTNm4lYWkvoUZBVnUmTONZX8pEvukrsZUnksNlcsadxnDgjlVz6yv3pOA3fir/Q9r1FrQjt26
cdMrrRGYbzFBKK5BYrmTsPeY2AC5XdKc7oE0WfaoXTmUvjWfkzU29Jv7JGZIMxoUrCpy4dgUnJxh
cgirHXJmblxmnvDQaHqN/HVWrO8Fx4LoEMueor+lojootj66K5+xHqPmuI3BvFVaysnNDQ3hFLXn
RfoWDWGVX9Q0xBdw6oSwq8N8NP4mlhpH8qaQ7Fv7asBRLtjtBbyYLLOaCoUFih2OrYDw6Bv8/hdD
fvJ+/toQ8kw6NzcaAf3YHJpcA3y+tiBpRoUthuUdDBnNbWmxAldSHRPX/VBJW0cAhG6u0aq1rd9n
JMQ2AofjK0kBnaQerHwwqGhHIiiIikCdx7uByaf7OGFz5fMoyVZiwhWU2Qk6awcHddLtdxaKn6GU
u3cjFQUsd69c9zdwpprxM8sUM2jHDsCfxoNjG/j2/4qPgi+Pl1gVXNh4l0dgMcHmV5rXkdc+nJ/z
mIsnXr9OYhaL8QTeRqcUXggGaeXjc7Sj8lPybQb+6mCHFXitJD/ql481fkFpTyCMq0Xyc/G473V5
1mpw0T0KiFC5aPV4Fq8GBgWug7olmOIO75OtxlbBQqhvVfFFjMs3n6womOHQ2M/zYy0H6q/GkUlG
UbjWcTbiBdbfuuay7DYfKvfdBVZoq1t7WVMuLhSv1AOHhaUC6phOEVhbodbTRNXlZho9Ii/yPJyN
9h4bUeOjTAULuoqpaNhb6ooE2R9sgf+1wUNk5lPcwXXw8UV6vDWfGfncVQX828RyFvTKQJif+8kO
upL466ctRlD1UVrJvomlNmXRJV5fETHO5lNlmIHOHExFixCvZBu2Yi41GRdrNggc76swsAvnCe8J
K1BzA1nosYZv6YjbrpPpcJ3i51t+AwJom58At9wXzbC6Yr98sfb7NHj6uljhKFfXMf4CWtg3DJWU
PaYnXdHZoLw0ESTniC6Uh85QD4t0B+oX9txv/c/QKhn1Wt/Ayi7kN2ROV8Lck1dQnkWhV77he203
3ibaumE58X1aED3Mjk7sSIaH2lKT1U8TmfvJysBxlz7sMx8oqqvszECoNnth/iApyaKpvw79cG3c
9nXiT+HA3c7C3qwHDvqAQ3K9su69nC0kZTweZEQca71fIEdhNDYTHehXJ9aQcCqzaOD7xP6u++2z
A+VmAa1gPAqcGSA+/ZP88LqP+2LYzJCiRS85l52MA75rQfrMCgTX9MdNIXZq/51McY0Clzh2KLiB
EQV3y2yqWy9guFBVHOe46ecmR9tMtH0CTCtcCfKlbrQqJo8BDpLav0fPfNpuG3Rehl0or1KikRJD
CwI5sYUCngZZSI5hl3d7zcBElErwUQ+tvos4uM9G3yzHoO6m1g6joGnweLiz03xzoNXa3qEJJARq
l9ClmFXP0S76b2EycLfBOMzodzbxvtKtGNIKI+hWkFWY0uBfz77EEavkOx98pUdevBZy+XlI/2ti
l6SLS1ijkmxUyWncgUOmIeL9effmbFXDbAU1qDvqAz/COGcNNUq1R+gO6/2m1gRbWWOETCrrbN1q
Bg8zunzmrS91J56+k4fisury1FQy84im/LvYl5IIJLxcFNowMAoQ6Re2L+d8aUuFoH3/PP24X/Mn
AT40Yzoggs2TSngGQAtoQJHZsQ2Q5r9TvopvceVXh4CRJX1DfnbSRQMbz2Kan0B73pSLAp/FiV4c
NZ2Ln1IpZTFtgwK9dTJeBx34Ufn3LTfBQmnIXigWdGNmSCHiaHrhnrT+mMGL00sHqNw3oyw9QRr4
0mkDVza4SdQfmAcFmvHlhbxziJUgj1xIbEBIj+Dp7lIlEi1zzVTx2oDZ/GMFvaagcLAzvI/Xm35f
4YaJ6MGznnHhAKopZ2grasgzdHSt7dzBaC5M33ENrIhz69/fFei0J84zH4HF0+FlomWDO9BYic3d
LsZB/wExzIZMCEZb3IesqFeAcQtq3dqDmXj/N8S8kzsX5BAoF6JPx48k5oukoyj0pHDK94qfNvCK
GT4c7FceB0Z9BCB1+ghhR5vuBRcDkkrtnh8ZzkK2w7NDskP3tfXJABhIrr6QMTBNi+LAZDtETcAw
Sf3fBgAGG5tfpBNSD0auLOk6tLv6NHPDkDr/m2NMWsz2Hs+4Pxjj9n5RRyvAwdbibt1/QV5Ymg1f
l0QdhWbz6YZHY5/Md0l3yBPFRhx8bN0qlF5zfLTXvUL+JsVnZjrEFTVY8c4WzCOzPOYJ0mwMFLsb
DW9hgvtOX5UrUIet7KUMMpers8CKY7hsKgA6sfhve5hQ2vJDr1WxETzLmwyk1tac4DvS+gr/ek74
eG8AaxWMcgL0nmPkI3te/Dojy0JQXTxo0vLFr0KFGEYTR2gmUVsUhYthhH9zkQqKe1wCoL1vbKmO
TJBaWDMP3wmzzFQNaEgMiHR4hodFMV114N9DXfpxGNdWP5/49Ia8zMy7KQ1ON4pd2pj6r9OMfO1D
BqfPAWHvDpBfK5b7xsRrwwSgXVEu9ciFjWq/UApbXypYSwDLtAuxufGSI4U+TYBNS9GDZf+HflpV
MuVwNGklt4LfU/TqBsRJRvchISECiN6PARRapxGcHyh7oJGAVvg0vQLVf2+BzVeIawNegezRqNAd
Oc7nHBuXL5prhGTGCLOyKzMB/pscb7QkVZvG8USGIjeWRMXvg3i/Dbm3TgVdlVbsSGagPhh6EDDO
AoLQHRaFp9ra6mg87RR4y9koWphJBDjEyn/LtWa3cALbyNzz3SILOXgxqxwa/+PqDCI0rFfkycZ2
J40ObfGlDCcK+ekDea1/O/KVyy8OCKju6eOqqV0vn2eZgC+gJaM1z7Er2D73aFBBfFgWCy5lpLYh
OFpsgXcyFZKI+LB+0NVsWszwQkeAoTA8z9bQ5BCWHtN7W3gc8y/4OcNH54bqhpscHbrkbaoqteHq
7CJpVGS4CN84iOHstmrcvZpqjbsh4zseD7evPRQfvJKs1zaUy+oiMqqHIW01/H/hnLwvnHbR1qPv
pi+Cq4PgBq0smyBjLuIKfDtymxRxtNwTNx7PyT1+ziteSc1+D2tYDRtUjzr46YJSb0Lkfeub+BRs
B7TpfvtUnTZjqOddqR/a4sOo2T8agpe0u6QQy3MkLXxXatJzwl8aY8OgW7lWPbhgP90wCnACiglG
+ycd+2G+SVeFNE8+jc7eN7qCr14Qs50cubFsuFMthu0F6yntacz0WYQC97lLcFQoIBl/Fqq03Toa
X5/wdUe/nRWlHYX4ap2sKX1c7ypttlvIhRrkk52IL3r9WwCi6sS8RjTdlEanTgA5RmqvEdJZ+nuF
a7X7Rgz66I/slg0/ebgmG+BwD3Gu4UmQw8nLjB8KzfSd7Zd7nymuDcZGL1xuFVPy1hFcS1HMnEnz
vlUE+NsENRSfSIUlnIzokSTj7vtnPa+oje/QiR1FnjVPwI5SeSwqseDs6TAD5I11+A6ab0H38vds
mTgssqyW+P2raq4LVtgy3BFEovE71bQM6A+liZFJNhAXfv+ejse4GWTcAIAW0fz3/FFn55191T0G
cN84qZBkgxz/B/CZ6SbiMewlDL3aecegnO2h6t3SUeQp0p6WPY0bTB7oUAP5cvAYaKNFWNOkUR4d
ML+2E6gxuCwbzuVsWaljULAVsxJ5cU6ZB/78exT46nKk9c3pt7KGJ9zAWl6XLKuiIFCv+15l+GMx
oyCUvEz6FVCFxCdxYHDDB7W4zo+m3kXAdFAsdErJrDyCPi09WaofUTOfbRtj/+TNEK6FZ7XcQCOA
ITsH25totY6+1jWz5+ZL4RhMDnZItZ9bVGXvxyQMlY0bvZeKdw9Xu3phbFdUd9ngsJgtSYECqmS0
A7Lj/u2OP+k5Q/HifRtgmUTvmGOgA/F1/bCZxIuXmdn2yQBw1vfhsjK2PzikEF9tS4cP5M3ozlQU
Bep/d629cWLhRsaoK19zhwkpy79WE/Awanox3IuIc5t4D1jbRNWvooNFIphU5g7fR3keI9dPTmMt
w7NRzcGyVg+NudMbXwlQ4A4DbnXFXwXhSZ7RGgi1PaUhHose32KusmJDXFajQ0efcNlsXzjbzrPa
mDxzSZRvp/Sal2nYWB4F3Daz9zSzNCn9L4H/f3hpJrsg48HqtYh2YRTgAhdyzg1mSDn/EKPI+aFW
37y5z+OCDjR9d0NSZX8dPFV7NrLQ3Xr3tbb1w8kU7NaWszmbf0okisj1cmUCzu3iPHG+4/K8tpjA
aPoXQxdFcWuQyOxsZM5J82bY91mfTffONKpQgCMhp7CbIn0ATb2VQcK7ca4uwxjHFFIe/LCTvynj
TNtFZDSN7hw4Bt1jsn6NE+H0fZVLNrkbALK0E9xC36t4vx5BjAhTOsfvbavYj03VTNa0KFHDO7Qh
R0tz52N5qX0beNiUrJ2zdLZPQB0owJyhV2qbfvwRlQm0X2PIiCnMXbs+tp9H/HlaF+0KpKgyFdL/
9J9oO/slvy8LKIg+6+17mojDvdtxfdlik006mydeI+885nIIV/BW2yqNwlCMAdglQXf0OoxwGzRQ
UDE1krwNvd+a5UqKuKGUPUwte1qGTdaJzb7XVZRPb++t+QMje2JXQx0tqf7GH7vGdWizKVMuJEz3
FFfdsNVTJqwdFZ6IFDvhqOT3E3KLfpn1PNOQ/qzYTJcPfHAjfEflZ2VMtDCGCtBXWlkIbz//4rBF
apb4dQse4886PGaFjRZjJqQBBufPngRsOsmrerPhIdc/7TwQezMQ2M9r0u4MI6C+YO2vFcpOYRjh
0IDLcePFZcCF8S9HG+5kp+PThi5XP91OVZuB4JPRntwNgeNONhHjhUsK/ww/HuUIjBEHQT/gYLq0
+WeiQTpbv52yQ5evimGTfN2dRy2iteqdVgyIsgeW3gm37V8qoi0FGPKvNOGz1XnVGoR8+G7es/Os
a3jLBvwJGuA+Eb8fCoBwN5uSBnNps8YbjFhAvluGFsgoI5W6VEcW+QNloEwU9XVKIUN0jx7jfsgF
PSESkaO8MSNdUQ+N8AY2vz/wsSC2lb4eEt+4t+0fK8sZ8CjLSX4DjVRZkLUGS57Bc1bd+W6WNMDW
VKqNXOTaAdut3LoaXeogpFv+5bWBtGZ4xNYI69stB1wLONgvWNxch8zvjrvR2G81xj4iSRgMiuD0
jn0rV+I0YDEgcng23UVSYro8BcwYTUjOmXV0mLOPoYGDgnB1qBL9OoZTrQbuqF6s9lZfI+ycOwqW
9Y6p2Ivk6s08uni75F0jD4S9HebdZwqeTEdjb+o/bjA1QUty5Zw7G2mjg2dDiCs/XuvHpvbQyBb3
tk/D7bhwrk/l6JcqYa94beMm+HGhu+oLyhDiSSNUjPX4OO3cU6RWTd+WIuSIjskTz5BhFAFdkzCg
EIbrQkbTkWKHZh06tUvK6RNWlPZcr9PkHkFwOmLwK8y5o9oP19N2bWmBU0URTVkQ/y0fm3xA6DjS
74zBZx50p0Rx0SVa5CtzsgSDB++vzb0fcJUIDitfvCmpSF++VW7BLX+zcXM4FUWPedNCPBwbHT3k
Fl3rnpLjl/vKkD4sj247zWHmM2I55KWRHPAsSxhyD4fUPtTaaCfjUwaRcZgCGnk4PxlOc2JgBqCT
vswLrKLhNM+/43BVav1OTVcEMiymMipufkgMHTrmHGUvPxORIN2P5hGrXgVPNTJk0uwNyPj5XxzU
1ZxSsCSSMmbRqZkIRNdqeSgaFRAUt6uWUZANxwcQXnTup9ph0TWXXcB10vPmWkxh8QOdVnJNebz1
MhUdlhdzdrEsVYnRwh+FC/NSOke31DTbJ/hA/2s8THoBoOWCtPTp1r/bUIKmlyZtMziDVk04fudA
nk+b9wJW329D1Q/e6RI7/PMrRMDGR75g8nmhwFRxTqSaimAbxuTyavuFlh42tnt/75xuB/dJneW4
M7ACLCASB28B+UAaiOblbrFVddlArSvnEkNdPXKa7YAJ5ZOwHzaLQYvzgCDrbcXI7iv4o4jFe8J+
nMKZhJB3HNREjSJ6k6Q+L1VSSPGfpqfk1N4tBNmEJleWw/OReADClD97ialAgbopM9dImvsjJpYt
tgNlSirF+8AR/cBhtXjpdLYxjYsXKo07Y5b1LBYmzQIWFhFME4rvkrnIpS1XT2M1IMWBZdJ7BAaj
ChKL2E+HDO3Q/Xj8CRPv8CBu89ZNolewUOD7NSPFORBDW+2dN4BqKzLBESi9yzN0GmS6YRpTJhgC
5naB4rAUc/MN36Whn9eoANI2lshO9kALreaCwpAcO6am/2E4Yda3JhR/9JjdivS3R5Agibv4QgEV
v/OVzU64bKX2lrQHDpSuCsPrFe5N01nsLrimp8cfhFKuTaVyZifkJYR2ebRcD4iUkLAM97U1EIpN
wc4erXkAoTTFGR0mNYoNuLi+qA+lDK28GyiAcjHtmiMfJIu58zlpLU1JDwa4F7TLIdeIExML3uvq
w6aJa0kM4HMleTiEUWqAuB8Sc0susEOb28RTyOPUwktXx6dAPq20PIF9f0f+8vIgl7SMd20GyNvJ
W5KxDHiE9QpEsWCLKdNYvVPZjPeqldqUJR4AVet/R5DlFuwTSG68+LFnxftL5DrnP6f4Yoy1CpYC
DgxRrKd4TvyKFy3WJhItdKqbfkXYOqFKHK8UobGaeEDu3MS9P6kc7CyTNhY8lFfRoU3+kOjW1Zau
+jUlNtwPt18/rqokPzRdcm12lm0hzPws54404ndCSjnGODKEXM6R57WDbtlUPDf79KlujWbXEdk4
lq1iDivKGKGHvo+Atd63SXKXHBjayhOIMf1kk7KdNDf1s66DIOfiwlqgnd2tMo0CXOMj7HFFvM1q
XWbHznK7Mud6jZ5OvO7CGfxk1Td+VMnYToC6omF93f/F+DW0cx7qqDbuReeMWty0NCqbzkDxoBgl
SGDn0w4/LD+M70jnDrlWijKVHNR6uLMKPVGthV8ZEyLXQJ1ftzHK/FAybO63Z9layE0VS/2iLGFD
M0DeHHI3a1U+TMTK7ykFhGerFCK6dHQ1mUTrnMusOPKLBvsGhW77IsJxQ+vbjLnZQC5W9MrXGEIp
pZoIxKGKH+i23HdTVS31ZGymjz4WzaoqtJhqbYOra0VpA/MQtamIR7YctT9O2LOtDvl+I+fI5y0S
KuTe7SkYyvuhwvBwFj+EoNnlMAyrVYpE5vAXeiNT757NkKywABKbdz21nxgaOaRmFF4lXutZ4Fz1
biTG9xc4Gx8p2nbpypC+TO17x+BHlRy2dKGwHy4IjTf45xsGwl19xSE1HWGg+AEOn1qnx0v2VLZZ
EuF+RciYrdyyM53YdkSzmGxcc8lvqGq9QxGaagXBwqxQ7IpUZU/in2stpohWv+P9ERbPomwn4dn0
FXEMiLrmbgQK6sXw+WekCfV2h50KjLXDZ6xB71uCxbQK+gbRG9a+cCxvLnO73YATnYuiQunbqWiH
uA9DgT6RCxoViiKftP7sj83epcmnOcnALDWMGOm+qQy6ZfDhHm7kDoCnZsPiSK7/QqbQZPE+wN1E
D8GaHKVfPfpH2i1ZkG2h78TLnhffPCuugHhi2cSvX9JrZmm44t0+nTfJ3laRxImclksCIjRfOkYz
tHrlhVEvJJN5H6XP5cfU6bnwr/SdJvo5Gx6lIjT/dUBJkALWrqZ7+LGEUqbCBTI4+PQWtqEnJDmB
+iAug31NvuD1WrU9kjb8hY1D4QQcWf+8W7gqJg04evg/Nht5wUQMwGdv2ob0Q3BQvPX/OE7gKPmk
tH+gxZmEMWIE8FkGnDvvuRyjPpT0aJjDWxx43Wk2bbrA6j+ipEspWiIx1S+VVzQirvksVXUfYFOC
mz22saHs7flP7f5CBtjZFT1MiErBHMAhhsXkoPCPwToOqGdNnX+RKDenXcdjeGCnWZSSQseDofh2
uRbSOoa9RTVa2YNpNwF6IfZNik+5XkIhrtEdTUMy/eeqhJeMbiU4gA5MTz3Zky2NowqreTaW56ud
AP5KAnmanXFtGCn41/pHoor3FakOrDoVExQGRIUrTiHNjUioW+rpCs0jFzGRaucwigygEtK91QG4
8Dq2nvhJqQabQUKHMRrqI8haux7c1feTmR1jZCBQGJ9pzDCD2ca+ej/2Y81WrhkfAVmD1HPHfHIh
VTdWNz+iAVqrjy2ZNyQ7IIJNja5uQJQu/ZPnYjhLTj76DvtpS8cJrtptdJmFXuoguQi74fwxdW0g
CseiErBg321zVlql49irBG0xfQJn4iJMcbrdqmhJLLLgRWiEvGnOCMVZw4/wllugSUT1h+3CEKru
Hvkk0ro7pGvLGfBxmYXyzLgvrLzjLlOTdfcJoNEDwd714KbaQCCdj5vFcs4jSXPCs/x3V6QqwLkz
zyOfBaRUhWt499Rk8fg0K8u/79plue/gd4g4FzBm6Ct52uurfkeRt8Fe14yARUuzXB7Rc/SggZVn
XwaE/k8F3upXkcgO1AOBeQGWsmHDCwByoq0B4gPAAcIcypjRumGeut0Hp2YXoeTHtGVdyCMiQw1p
TdsU/bDED8MFE3WV0Wax1rKM5aFuCHyiPopryZYlkeymK0+3Y6EKcQTAfM7xmf634drd8CtfqXxk
3khg+ExeknMuo98HJWsZeskXsg9ah9b4h+za8r2aSuhXizd08tMVFv8ZyNUpgEkvjjR+zokjmLBu
9jbGhomcBuSgIheTmp7jNn569ASfINfqDeS+qlNQfP03493l0XP49tWtn2xvo0qyZ/mfM/9vE9+g
HogpXO/Jixc0uNHcCsfCet67MkTw199E55dLEYtRHGux05IU8OzykLnAwiKX0ftE/koqP1CHOiOY
YwC/HblgYUm1QbwRnZ322mrbLitDnLXkHZe4JGiHCTFI7OHhPqqvYEdAnxgatL/xWC1kqeCZLzqs
7R2+P9Jl+wTU2H1k+6bjSs8mNKcStTliSh9DjUVcRYLGdrrq1zDlDbAUO1JPvR6WtwS3CwJy3ET7
3xNqPgz7NYqemry7JX4Trltv+SP+elKxEIOSkhy54kkx0yUcI7k/1LVKJxT2W+8eMSrgwhbIUcsv
Qyx84/DO04ih+Y81kHGMTe6iJkYJaWqJZFZQ/YJo7WwLjQUFYB4M/5oMeSxN6fqPspkfJXDEC1Di
yvi/WAqeqhhjxUs0lHbUDT4HreJLuXDqVB5fZ4W/iWx7MOCMzrFeEXJY4P20sGeGIU1s3hIrta3q
WCIz3ooocoaGVLNRTg+KWd27xsQXS6dhibw+2t0x5lT30gQV8H/KCOcnSaDAG5HpZx3wfsPL+aKS
w96b3bp/SRq9y+8sSw96Kzt0dMRTANRmMDlEoFDDdE2zZE44xD1dv4rPs7N5PksOUR8EXvcSXVxR
9gVFsTCdwvCUk+72Tmo/cJ+b3dORSLSkqiFesW3vcld0phA0oBDWBB3GyHDlj9eLas5rNmL3EK7S
/zYf4awVgSQV4OSltEiKq+uiPrtBmPKoFot6luP5mQaPyJlLfsmFwCNCp4hh3eBWuP8hIKZNjRe0
uk6YHSPhJNqd9VX286qvzzTxzTB7ll0NqBEVusqhhmWfK60jOyb9ZTraoyJe2p5vtdCWAIhv5qBp
8iOyfNxRz4sFerK6V9zq3z7c/vp9pQxJYSJn8+KT9DF3maUG6yypoHjGbL8MV1FEL8FrqrAaFaS4
F604my940T1+XmHwkgxj0GB8JKx2SZfZ3ISn7G9TrYLT6H4xcV3ser0jApfdayiFrjLxV1r7XZ1y
dvQ4b0lJ/EvDboUUOO+aDemQr4EBziGIZ4m1SUeZShH/4+YMF60BZFOInTxaKbFrX+P+6lg9o2Ki
2x2eQ9PuKsJqV8h2EYD0Pd+F7uyRk9NlGVG8h4TJ5KB/w9IyEqYP1zWppXX3tHEfE7awjXIYhKjA
wlfvw5C23SnoRA9bzVrTwXtWy1uXC7UEqEqFRGrDSO6XZ3lSR5A62OhSoXUnO5gJ27cf1ndgzQ4K
1IcDCPNxPN9WZWF93+4s8HyTILVvxw224/tEOPZhXLKBwiZwAVGr/mLgCvP96gCAWdq7nJicqVRm
9qZTxZodJVVpkHEng+6FZ8hpYHrjeGABBNvLI8Dq0SD0K5BHqtIre6MEjXhS86KxocK2Z0a+i8He
YeGmDHsQeseON6blRZNhrk8otonXSdYUUYenbPnpR0tpUHtw0PNbUBDrPseXN7iGB6NcvIiGQiPT
lQLhEj1/javDLVvR/TCLWbreaUuXcCfC7r0I2pWizl+R6FelLEj2115jRF8o4IcronpjdXJTZsYg
HBBxaXKeH/JDFuoL4tah5U7R+Lf1cOlzjjjaa5MOFLCi57euYd56Zoc0rI5AEaQ75f7xZ+U3FG2Q
2N/Xs2T0a4QjwMF59iEEAtnO6Xh6taXh9/raZDMYaEPZ5HNVBfpvh8dc+hwhxQ+WI/B5tW+fHwyJ
AQHP/r/9LhThOylYR6o4AVIH045+0ur5zSP0CzMGG/WxAVox6GGzwa2I4oNRrubo0O37VVyQPxIL
f1Ltj/Kw3m6ru8d3ogEcuKJiY/l2KHs7Z2UlpV3G6KQcIpcRXZYTMIX7jzGvrMcdm/HhRnthHJe/
iVa4jft/F2gpdznr4izWpY1KifspLY85AzjEzd85HFHwa8itsW9Dva4+VNH6Y9wkof7SXBdzw8xr
fM5i1Qo7DhFgY4tJOT1dWJDoF3ED614rgGmx8aqweW9wY9T1IJWYEk2xu8EAM8XJxHUDH4g1lATR
boVZ+RajXdD6bEobSM5+fSTruzmsqxpOfx1wonXmr+z34zwg+i/ffJUurcKwUVQ4nBD67Vc1wBup
+82bnlRRCQTZCh4i5KBAB/NLXjIXSEcIjqfuxFoWaVJaaJcttn7+09NX4YVD7JgOSXLmHfDdkA4n
rM1Zp9wUL4FoN5AOkuoxyKUk837ASDS1biLJd9BPVKEjWddsSNgIWeCEg4nJ96L0p1eW8WLCK7Dt
/lo1PpRcDsS90pg+7K4o3HrNq7A4+gqhUF8Wbi/430HiQ4XXX3oj4pF+JQxEfOLzfM5xu2H5rx7Q
MYxr9Mv5UOtnSc0Vrg1hIy1hoiBi7XrY2qVy93KRzYtZEqwarjRXiS07i4D8vAK7bSCmTXYtgVde
fHgwCdV5EXzgsAo5I6Jhuvy9VGNEDzaDuITMkxUZX40I192PAel0ft0GV+Pn2uhywG0EgK/z6vI7
uaV2KoFIXFLGBtL7UAjZYEM5PxxJiW0O4TtUa/YAgiOw7r340o2hKtLe8ZevC2LymnLjVym6pai8
GOnu/ufUcvBWKb1dTq/Cy5CLNp0X+WamYAbCIPKQX75oF0+BGcWq3YNgIrBUOHFAZ86pQLOdxkXn
Eo9ZI2Gp0IFSEkmVxXrpf65vSK6UEJl9/Y2DPHkMX8bwzglE/ifhymvAd6lJixDdgmLHhW8B+Hc0
201uOWlfiT/cdrxEhxnanYjqnWXvqa9/uT0a+aIzuQcCww1nE7cGDI2zIEp/Y3irEZC5Fy4OGi7u
vqBshkUc9EFAjuK+6gS7bCclu8VyvA5pFFCjjRxQd4+6dg4tgXlXW2c4tNHrDCR1WAm+EQgC4DmA
+/ahQIn8mMOpBtu441vgmV4NhtaIvaAvGQILcKa8gXuU8jW8AuF8iVrV5X1s+R+pBJhvK0/awhvd
143NipBiRMa8Hr7egMWL57VSERp3hmK3ZVlIttTHITLNcfVUNC2yfoS6/heSVh9RssxcxffkJZmS
/AALXDQwPDeFTKk/QXw0RxpYD5qVeb+SNrIaNoVWtBJ3Jnu4ussv2ayCarA4pmsopNWGDkJ/4ftl
7O3rZD5XsEif+dg0KZH92D5liXAj83NUEyjLvP+qXJ9rLshA6uPd9sWuCtcXwwbyONPnRSzJYqfk
YiEXXKhTUveqAyTImv/wUp8ujXjVNMaHR1nd0U9lQoUDNyUuRIEOy1C40wf22/bU0yQor1zFMuY5
t5UnK5mUQQb/PcnEYG2/TxXhf6ee1Z2xTZEbioAm84ZEyRFenV+wute4J4HICgEL/GEUroeUrB7V
aYVKfbGkyfYMd5sZFuvLsLMxhFeEnM+Wa5htjzXjo61ksq/G1G1OYFP4c62BhnKbBwHa2RomhcyY
yvnIjoLussEgrgkMB8dPh6Hp0J22tezlK83mVcouzuQ6WGFqxq0jl/4nm7OlOK7TXJgnRC8ErQ2c
wHWH2KHmLGV202B1zbLXf/17J49Fmnf7w63ZhP7T6NIwS4F9qFIZx4T5mvTRKd/pno3fBM17hXPb
kcI4Unj6uglHW64ilCQR21OiH4VV2gduMpmkQzgwzjJXuQV07Z+l9FUcuDOgpQ62bO2ch15YEnDg
echWJX+tOGdn4Nm589YfVZcWxb/J9Z0KV9Vhii58uoRNs9yleta5tN47CxXAv4Vp5a5Gvn5gVWOa
I+c5rrGbqHXz7OwguqIiq9WhRsdfXnwyIZt6+eZkR0Zb0sS+5xLrKmecNVt8pgxKpWQ0ljqM8cEJ
mYmQi3zW49q4IwPZoH9NrE3t8pjiMtZRMAa6Ib+R4r/Z+I0zA9ysN83yHvhNlqS4ZOn2tfQzmtNA
JgzBrbiT4ZejeGxRptwJJNKRQGSZr/+XQpUfr8AxEQmm9rmEUSaSTDH7VvgmkYyNFItFP76MB2bk
hdsg04PamZYXvicLDY/g73PH1x/+bbow5hLD/haOpXgOXhF0y+x47rHEuE3rm/dIgDFhBvnF2pqU
ZfMQf0cJ+hl+XC+EiPtbESejtD34BAMsr3oIz12GS1CvwFeZ+e58y//zAXBFQsQscktov1B/ZgMC
x2mGla+5OXJJPd0NPi6wA3aISnxTH8XsahgLahVbqnaThabIpGinOV8RRkbBiwlYDeQkbBYaJ/t0
fk6BdBiwMeFypQzz4rvgVBatfPuToDw33QiUetmpx5BvNiR+efQfPBf4UahtcGfeanlu3MStcwAV
zKw/lIB/AAviYvwASDhFN3hHrF7ntw7ZIQ1CcOxWQ9FgYJZYPA8vLC24kno/fzvDNCAL1R8h7/1I
sU4L8QvgAbUC4Fk47tvp1V0jnmoYTx0ic/n6Y1J0o98ZhIeAlBN412OLQtq1+eGMR9Rcy/7fQBzU
vWlg7y5Pqozd7B6KlsTaxRm6wUArsJnnDIWimRkfLLdBGq8SGn/iycE1SM4y8J5NXZQrBvNjAR4T
DQg59rcsPiBfXkTYGkOxIGpJCOT+tEUOXVQpTnpiJLcmZmjew8blbAchHASOWQxEokiAdGmlL7Lm
vHX68zzqJBgCAlj32RWUtD5nIh3iozGM9dsVoUXTOK0x++Lk/QreYQcMbcp5QsdsYfOCCQFHUbdV
vpL0ybCy8BHC8jHbwuo1HFhZH5GKDXR0jGXRtRL98apOWyZQKzSZKkug+u9LMTu9lukNxCjTy/TL
x1Cjt9KuDuMDDgPFpzS49CtpcTh1oXRxE34lmfRhZ4UAzNLoOl8pb0DmG4eYUWSgE0RfbdEcQn5F
litTMqsZXXZuBXXIBmzFeMK47O3dTz/Yoxu0froBy6nqEt8rp4gVfJEweaeQudWy8dQfwAcs4Veq
AwzuSeInV6XKgjUvJwNVjFfq2nd8ejhAPtRQhidH4DnsJf2jdmz7DJM+kMxlmkkquNbbbUpPPbsW
o3v7S9jVWcX+MQQDs08VGEuN/GWkC3zqC4+lU1YJ3Ahs/mM1pPqNJ/td/iLVo22C0OYlwvQoo/8T
tXc8d/g0kJAY19uu+IBhDhEkkmgZfcAOX+yvI30WGQckp4+T+WAig432n5cR1MbpVqb/KrXVDYlX
9Zg3M3yGFo7JUcV+rmz/dQqO4Mta5Qy49UgM6VolJb15bdzqPk5+MjOCs/QiXg8/Y37iPnVa674e
SHxGlIHvaaCTnAkE2QdpvlDDTBprT4Qd9dK3THTVTcpuInAVV0WEnchJ6IMWHMbRryNA0JAkYdzR
hZ1DDEYw7C9ZS+pLwXIsnSZmk9PVRwcs3nFJik3SrQdacxJHHX6u1QO5hIqZajVPEqbKl4eYl0iP
mSF5U2Sx6ZvszhundQGGg0UFmgXXK2F5Yd8YDRc+RnOAhGmXYGKyWJRDbpwvOyaAxUegl5nsL5lT
RLO7pwkyyyaNK0xgF18TiPcNpaCV9n1FwJ6HtDoe7roqkEZHchIN87+G9gdJBpkF+8oZZHxdZBF0
6RAmF3rIhRzS6MzhKPAyYmfoB3BRP0ZPkgvxTrQLDh9m3rQwCmc3a4OmoGVLQTU0CfQwAc8u3N3u
uRiArBeh4Fur2FOjdSuQCBupf3uDfod2k9wUPPk1eOaV9nGKqJkUiOgnhpxUboQZASu5LmE6P312
3hLjJu4G8Q9AtC1w891e1nI5SCZyLOG4FKfjP1j1Bor9bmJHy7sE9LVBSP61E9aIcLFVu3SzTFIB
Bq3lf8ahqKDl/edpLVTYy/WnMfztwE8Ds8/k5QD2hADjzm2jnfRqdX0hz+yXycy2SSReRZ4XsvFY
4tt+tFaBbugj2dGjpKOeUSf4rgqu0snxfVz0v9WlRN6LXpKs+Ze37D8fAxnkDRAqq00XBx9yFizg
CVCdBQqNR7o0j8z40UJRFhLWx68qMEqlTIxeb53P4UVSRrkzHwSP2x1OmP5UjFPa95qOmGc2UeIt
IGjdHNGp+iXVS7tRn1Zz9J9TIXazrY4Y0p2gtRGqguIMGuJ8miiYQSI2fq4Pp74uRRED1ETCA/+r
vtQo981d++xwx83mL4yvo3JCJ+dxU25iuxI5Z3AZ6DqwAOJAWK0Aa8NctSLdJIXnURVnJFDD84rC
1GnWm0zh3enMsmokrfaZTqEwen+JtU5xWd3WpCzhnngks6m+nOObiajYpLTBuLo5RLc9APCQqWzv
0AkaB5bE0H/ZpuJ909b2rSe/2drJkRUUhm4Q/sU1G1HXFaotV78gA07N5yXgf2Ru0gXqenWN5XRJ
FEaDiRA32kxRmENeKME9VDI5WAQrK3C0OSRqiUqAZffUHnhJnsV7EYO9k1Iw458ngvf3yZjQqwSK
kkL2U6hM1uDUdvWve8LFicW/9SNpjauo2YlGzDIap30dzpoD1GQAxhjbHV1C05j+fmdgatNG5AIb
U8sq1DgAf3LxbSsXJeUe/cQsyJpdN8EntnwrYzSsj/aM5o9kSrxUPyZO9/gSXS976vuYxd9H7XuK
ff5FFr8wbmBN0zCZBv2T9B0s5M7W4pCDa5M8s+gumPM+ga3OokuOWU9cr6xQMzvfMxuq8zK/qCXk
q0A82dMO7f4ZIw1IwVz2FJoGH21kUymtDP6tJQgCG3Y38qru6OzzfaBnSg3C+l3vt0VtOPDYZuNZ
veH4YjQsXzPsgIO6rZ/vBa5hgf9CxT75Y9ZnVoFLWwxzD83zuMtuKVO/F/qttuiF9pwybTlDey4x
FCiXIO4I4ZK2GC79IhG6VloIRIY+v0onWuj0wqGAtBkxOPM5aVeKPkV9ZI0wuwBEcp8mFrexT4GQ
ea6BB8PwDZgjXOln3/pU7yaZmRlxDx1yN5iApqgHBr0fQwiQY5K5om9AEuha39ppwToxMsxICpr4
7fRULgqI1q553Pn2QdC23b5t1TrrFMA13owZb8KzzSJlNvyM+mR9M53zHYg9b53QQuClhSM5gP1m
9yXIUR74LnyVtcme3QR2NkCDq9tMBHomuGvX7g8FWuTACxi3uHAsIR6/1gSuWhOMB9YgHb6F+hxy
vCZjBhD3X8N7BDLDdYsLBEWuJIyYuGbFBQHqmnjz04z1rYuEdSsygj/PNx8ShGtSFHIAabjdrz8o
fopGBujdUjzOVlTpImVy+Pty3WI4eyQnmAf0WqhwqpnvGPgUqoSubgy8ICpjRaWRe7y7jtqGk4xH
Ze5Ahx+yrg5u9xUo3YPi2CDVBVE1gq82R2WkeJb5xEl4XUYNpGU8XMIkCevw953tEUMR+FZM5Uro
6KL9gA+Z9J8sEzj6JjJsl40Tw95r83H/665hpNAklKSOe+XkZbOKWZWvG3Ls8zz7CUCk68G7Qn63
OV/kJg92ox2ilrcXuNZPLe5Sg/yIru0UtFrJUciKf21aorZeGl0oGkp52nrmjn2EwS4aA6P0NCl0
pBZtUDWOoPkXk7yaVd/f3hG5SInDq9j8j2Wt00eh1wqROC8L1VSJQ19ndiWgvV86KXv6w+UFg3mX
8pfuiPiiJBo8T0VLKV+32mIwCIayS8QbrfWDR4Sqt9k+9JIeVYtZnbqJ/X6FZwoXI06V3ZeLmz7v
D45tZVGSjMp5xxNpo9DNsh8Wg6SSjXYb0OzQAf23MCkzLGTGs7I6JnJ6hweM8Sl5BZBk68YoGjGo
bWEooxjqKgo0hDkz++h+fhJpts8vsKePAkyUg2o0XwT6DSj83lWgsJnNQcTDe1isRQ6zoreTyFzC
rralOkjlrWSyoRo9BB+khT8YtOQ7Lctsx++3LEhrUc6yvW7L5ltvq3468QLOhSpsbqOynf2DQwUN
L1QJ1bp96rvPEZFbignnSZvSagS7kH8MPjlLq5INp6DSOUeXFJGoMRWMInrbnUfUin0HKuifQLAm
YKDGgvedz7YTMMaAqfDiEdHD1uxIY2aJ8vCkwC2KT4NBO+CnY3B4KGR5nuYRsVneDRAvJb5e+Z3e
ZqpdtMALHeHCdXSkl7meQ+9ekQIC4KKMdMv2KyVvxhM29tocewhHcocsZn1JBjXtvfr0lVLEKryz
E/zdOAp2maekXjZz2OXqlPuc5ks41imCGFD4YBmiXkiZsDMmf8qrCh8GWigdRl6QaYgqF+i0zgqo
mfk+s91Egdr1jJNP1AnwfVvn63rHb0GRR4qJREB8VB3s6GG6h140OR0m04TTFQRd35ozGTvCS7wC
hutwM7qNsB8u/gz2fjUUo3VXQ2sfooyw5UGq7+/y4kl/3yMJzN0TreOIZjUNyPgVMVVN4CRVZTgD
cq97JS2wlnK6jrtrN1QSlAFavqfvUDCj/f2TOS4wl0lotLjSb8Le/Z4V/Pm6M5dUgaDFwXPkHP9B
2ejRXcIzbdiLdb1c5sgQC/v6uS0QGK1R7ciQnMesL6RJH+W3i3WNjkthgWZnMtMoGr3gIMedpwiF
+LGgq5eE7ZJBbVr4uD2guzxhWW/ZH6x+a2k0dgtnhChzKYNV1ROfw/JAxAaLP++uyEeGbCZ0z8qd
xLnRxeGP9yXPagQ6VfPEHk3EjQAyXC6Ixo06IdnGWjbzfbavveD9V//HM6569Z3jJaxj3u7CNocg
09N/ZHTQclsncIENgjqaMFxvayEIVclYwXiIT+XwH6l3kuJlvL9jc1nLMo08b9AIEaqQHyQd9l7h
FcSWIklyOdJ5Il7fSNWJWzpM9ifn4mm9U6NRDDL1GMPYTkt1njVi9+iJhqMh9SvhbqhWgxax/WGP
F3Z8ghZM9zwFWDijObcuyoaF7TrRlJPMPPq4WF/wurNICfdTaVCI3WpPAuPSdqM8iuf78Fy9xei0
R1fVz8Vr/bYvacjXVchBWr1ngcGQj/FO1GokdOpLEMxoP5LDp8eLie0wuKp1K1C7dqRemijzr1CP
ZL++9BveakWREK7BR3X31gzFF0HBZ3bQp++OgysdG1eePnEmucIH2v5HDiHrposbvyJ74IteilqM
nAtLLpefYQTN0Koh7zX88tmryQ9yDt2pWClbP2T//0Upeun19hXvR9KLUkEYtFRqooMjPn/kjx32
NzHb51jWb21D5mQXRytpIuozXChxF+BJK8TrvxEwDLGfeW2EnXPR/zXkdb2GJMxam3nbPQRrWi2n
QtE+5GnIyYJNNiaaVhkK9AAOA+DO8iIlpHLLCgMwYOcT9ddvI/ZxbhPjY++qSlSP3Cbw0ZgRD378
Wq740p4AnvKkbI5m9jKBMdI7Wqqe3MlXYJI4wk7WUInxIIzGXp1MN8twozebMLQ5+d0EYdhY81pR
aLuLOJHYNVt6fbgVogZ3jlihLFi/SH2uZ82AafZc4i1GpjptIIcdJFx8uJlrmlQJI/wl347/w+7Y
y8PZYW6BB+/QW1IyD262IVIYX7j+22dpvL/7bbTUPf12iqaIgZXe9rg4Itm7WhMeQuh4Fxjg2YZj
o1EPI3126s7JmNoTU9x842x/qIi/p8zvDZC7YSv+CTPfVz01nDKsDKTr3jaFBFU/H67S1puRQXtu
CqrE5AeDOW3U0XF8+piF0cGIG8dZttQ69R+aCxEuuzYHjgLC9Du7oD/aBurcsjg6J0PEWSCAcgcI
C2CxIHu1zCld/SrzPDa+PDSrsgv4KQzEB10nynOq6yArEVWvL4KxDInj1SeSuw5rZ7aLtZ27N6O/
ekRHCmCtFHrAOJnrhcxygMt+IWifSOK4xMJsq0r1VYElrkiWGB/dZlebaTdkjIpnTCup/x26CFie
pXeBJKFYqgJfuP9AyPKfao3bMffhgTLakYuhV3e/j70Hu4N0DvLNnHnNiobPAUG18goi406XsyPF
omfaVTLbYWCEXVLMH9Ajt94DVAi9D80xM5eqsenhIAE3pa/PGz1ylWodGM2QBDkt7soe+DXUxBgU
qOXJXO5FtE/R7hwWuuSGHzPkS3UEWNvZBTEcwfpeWLQFZV6y2HY+SHB8pi98ypWDj+e6lFmwX359
AinGcPtdVrGQGTiJrT2+CG39+oCHzYRgeBWQulSCB0iCnM7Rft6aSLEZDEyj+0I8NNW2MhLxGp7k
cop/7jPusW1ePap2MUPlJ2mKUvPSvfe2vcKt2NSwmQlyHelRpylL1ex43P0oGUeZA1jd9q5H68OM
SMTbNgTA6X5ccxOzQ2OHKVQL6YqZ8g8xsJG158FB/OWNP1vBTBG3XLycebMblH/MaJkBi2hV2QAH
wtrJ6o3FtloOqIz9TSlW5BEmjKg0AtnHzJt5Uo0PWb7sueO4kOmKRiJGlgnAbLS2MT2JsHvI6uwY
zlkOMJJzIOuFnhmYKWPc3u/cSflYlQ69loa3DnrxO5Ltlr98e8hF4bJHfko7izyj1oxonYMxPHbj
PW8RucQmDRD6NlTYc/IBU8/BKnCSagrrMWd3hj4LJFRh8Ga/w3ixstRAOXfvTIl2g7rBVJd4V0Lh
V7LatO9C+r6rxmkkyFdF4un9H+bOhVJ1ej+DbY2B8W7fw4/lj8jw12N1y9kysXyaisYn7JABwBAN
3gImbEkNo6tZJDLdFb2fTN92WEOC23xDAN0UbP/cf1g4ix/mBKDinABY4rJAYmPLk7E8bKrN+c/z
R0GUluVm0EJXOp9K5VkTgw4siU/POwuQQQCIs71sE+HQ4UwAgyqDJlQlJ//SMkK6exl7DlwrfApb
1di44yr67Co5h8ExvYKYYFz6tPU73FZ7tk9UAEM/InwppfbK6BDaIS5+dKrJ+waZ4/fHGTLZCz9b
5eg5gHmBdd9qI776EXhx6hVp61mp2bGGczLULyN0+RXxuZ/KFesAoTymDMvKUhWdek/JkK4PToBG
keWHy0cJg8seLizUwwziaQHarU/dyHvppG+6wi7n1E5h5MQ8IDHCN9mWtryA5Ha37aFKEPZ0adbc
H3y/MLkdQjc5vPPSfI33CF54fja/lsIt/5TrkNmxbuXmX3Jy0gSEYPTvepaKKXdh2Vdb0exVYnt4
Elky9nGVYfL0d4GOEJSxHjNOCVEEzwiZ4GkRy5Li5m4xU5m98oAvPS4K9lug9fm0t7waUPLf8Sgj
Z20irN4bBK6HSN4amIyMbIYfU7nkeHrVnPcptgcqcaB3694A0ErUhbDyuF+6eeMqIRmqtGe3hc+Z
M5dcKrsaUMGrOc5pbZgck88IqYUAQqkUs4382Bty35MaV599SfPciaxp3ajuUI7CjcB3U3MPXNtK
dCS8Uj+7/tQSDnxbX5Q0mhMp1BszFkFmsEZE+Ej72GlULDwhguyqUrqYNK288RzKMdAq8HQO8bgH
mwBjRSRaRWcz44H1gj0iCVUdXbY/WtjF7FL17D2YPSOeoG/uXR6PmWGFOca6+9Du1cF7KPmyFqTL
IX9bC7gHYrUMuXHvQV6YvCXJzPAr/6t01GMnJTvFSS5b5u2GHo+mulT/YOgoHYy0iqmtI08BQxG0
gtX8ABXOLz5xOyMi873BWjD53hHmUWcYBxBySfrf8NWZi03mnRsjpn5m51E0vHRYsVIjQojvDO/B
vCtijITKpzrQ4oRC+ZGE/uI9nYZVRMz6A8Lu7fa5HzWPJzGE4exjPeO0cm+2eEHZRhDdzz8S4OXE
wqOYwuvMEGx4ZG9EeaY2GVEwScu2j48+tasiK/xHnYziH5iGCiGaSuiflnudSLSSrR2vPJJwA31w
8iAvFp+QsU4Tggj040mmx26SnVOsTNZexrcrU2U7HkKaP6sp4+peEkzt+HpB6KSmDgfgz/1MrmDN
agk8/DsllTf1z+3M4yEQEaRbnwGq59vCK3G6ixAEdrGk3kh5EXKWEQmjR71O8azNajYDdyZAFcZE
lrALKKfgrKYQi9bqHV27tb4sdPl/cOxrjJ+41sS+ISDr5PjNcQrzyeU1TA0NtR20nqJvjPtRakbj
QiMwjC2tsu8VAY5EisxhqljpVSEwQ4imGL80fgrB0yGJ41J3x7MOZPEXLdnfajsGLhvBmii6Lxjy
c96vkO+iDcWvpVcD9ubM/UuPwfup9jow+/sQ39YOslpV1FASeRe6p7skyDisWnmqgSVnDy5ptUVk
1CPTU7yRiq4udL5MMY8wL8RolgbmEiURD+7f6Ux/fIAG0E6Hm294V0eeqP+MyLkBAuN+X8lAE06G
imV891D/KbuzLbIiKPkw9hEc6EFhP7ZMYaFoIYA2rqgNQPCpTY2aMAc/t9rlVM9HNIw5vV9G8OoN
5UPL9G2JqRmc97BIe3DMN8SXJxLuHGt7PSwCjj2qjzsM1FzC3HtRD/Zhv5RxzxqClFM08dk+m6P7
5VOW12i36o6mHYIiU2iwSO9OAmoYhANPN3ie37kg4PREOQVyKz/Fh8gF/I2DGxbak68IOLQO2H+l
zxuPp4GdffTyfFNdIHzrKXn4zCQ8LTinLVnWo8K96ntdHDTWLNnUl/Zr21RQLyKxBRUTjS1R5lnj
WN9gXlEDiqOjzMqb5cHAaHrVFzgPTx9Q3ix5ZMUD59WdQIKhjcTMmmrtDlWje0JWrShGzY59Raqk
4VPHXMEygfYdFdepHzYDNk8qQCTKpE1/9JP5CUk1ZaOWOPLn8Q5vl1ajENO6KFELYO9RdUB18OuW
IcVno+w5j52izaBiyDO2hQ2UE1CN9BiuFX8B9kzMOxGk+mnWFXsbYGNzgeMs3ihG0sxNJhFzx2Aw
pKE91z5oiQhdSIu/RU6z/MNDsKoix5al/cIfykrV2jP0aLwpcFGHSuhqv74/E0sP5MSZ8IkW02px
phw4i3r95mjbyla92gPq6xpfnSnmsduqwxwHRSJUg88b4ilGUn7WDLVn3jNuofmaQK1T36qwx7ta
rE6g/MKEV8dpuWeqAqrk9X/KyAsla1nMbqvTdilRXqtIjOgCKUX3I5wBZibqj6s8H/P6gDiiysbF
zbqXtNSKyCuxqyMOIImRIrLfyfRR/uEwbH3jy+wd30AGSQQxbm0tPUYu4zbnO7PPs0gHjCzAVic0
KbKdAj1vV+NTNC6MrwIIvjrzeFArEAmIwZJEshxuemkovJxSJA8/oJDvJQQJmgUjRd56ZEKepYSx
jCm66XgNSLBv7ZrCM3mEXXMQO+8QIoW+6gXv4tAvvpy12YnWhQSHMk/bEHB+v/6mWxrgpofMkNO4
o8qLnHKltCmnum2TfHqKAWwPwmmxM47wxHPiyNUv6pMb683XB1UGuBp8j+G4X2WtmZBC5qTivKyz
pu0v9+AD9eE7dxpTg2z3A4I6dlCHC5GUkVLby698D91XtnVeGAGELyx+lnTu126HXMedds4HeF1B
D3rLUPHOMyiS/c6tNepkDONI/V9K1/WGtzxRQd5UGmYvrIT7fA5BrPSeyDabVUiD2/pZKDMHsbJq
VD6j6LVPtvKDNJF5Xx1q+Sr7Wc+KCghPxxurRJBxIvHK1UhzJkZoTChdh0e9hrSDZOX2VmgtFHla
qr8UBtEuVdPaCzuPntb14FyFrcX/GgP8obBDjraLUz1Q71EyJZs0LaBovv32uSMzGEfCqSV7rLOb
4/PVSNk0NCo8yvTNM5KIBlfebuFOkDGQ0VxCPG/wyHNQasyBobpB9DlzjzO5ZqfvsthIFUOEZ8Mu
W1GHRj1hxsNVErdVgrgl+cpsZ0mNnUm3xeasGO3VdqFu0YkB+M9UKpSMW6IsUBOWEOJcZBzS3Enc
zddXMIbFmopMS1QMpsDJzurc76rk/Cx5XMzuf8W0EmfOLarEMffDu/M4F26qYlyPgoaBwmrLg3J0
ZWtEaPpAnpyM+IGJ6mu83Gz9THBI/IUESmj6qf28SAjwoLVxACF+ykBcDNrXBG0XPR7gymQspxPW
eZYlPbmgHyWOL1jAIsw7lm9O7cV0Si3mNIxxMLZR4kS4nSoA2j5ZgewDC41bNEv7kXmWH9YtEnKq
hmaBk2pAuTOF7q0PgI/FK6FRJI90drC80SUzFpVTyqZWFFBsPUZ3CzqCNe4syzYMk7WJ3/q/3XfF
X8FGgTAqlr5+i++dRG02Wpfhtgy3ihKlxEBXGMC8otT3ntnBohBpN9Fk5KBt6c5qph6s3HS2Hc1O
oDHchvE5tW19cxNh5OPLg5Qnaw91qfzT0fEvnGLX/MafVEaQ543VTouImpTCmGi9u/V2OmpMqwwT
CxZkvLcuJQbPLvjIb99hXpNj/7NLi2cR+3LCwrh+EeAfx7k8Gqf5v349GKwwEdlPHKWzUfnvrESl
knjz0kwQ12fPzljC7xdfEoEy5GQxdmRjs0O7dVX1wKqKO9lEA2y/MgPGjTFCIs8IURu5/fw09fMD
vmqVnRTJvtr0cqY43dbtFRrqf8PbJdd3K8B6/OZ+XDamOnQxfukvaNG1MksE1otZZfiTnTNzNnGK
/V1n+BCZbPAO34EcsAUvtu97O7cNrs+DmhmzFxJqTWw+lkykAvWtnTE6Py/5FtA2i1W5IkiuR4h3
E6fbWc2VFu9xt5WwJ4rm4Lw2cKBEkm+xyHGoY/cMxUJmFiy1D4AboNd+6BgS7mucj6XRzRgip8E8
DzER/XaoN0Worf2OUPmTXpgorUIGcBLrRDUqDeatQAa3jtgvj9dyjTncdsp9YFPiFSji8dsksKg8
Bxx1qVz/zmJO5cI5ZDbvUuD6RzEdpSOt6+GQMx7GX42WdtnKgxLUuIoDMVbaeDuzthkDt4VAnSpU
n7kqKyVlnqcdSqe7SwtNbf7o1O9NnArBiB3Ws3xJr4Pj6a/+3VdtQCcAGzeownIVmIX5pZGvN/Ac
nE8USFZYGznDgQFeyWAwo8bS7RG0JRjmQsz+sLbFlDy8whlAI+lua0lqsY9ZQFDqHlLhujRO/ZxI
Gyb34x4gnrbQV/lUW7n083rgK8JocLXBc779wFWm6C7784AJyQApeabRKL6EpT8qUZ5CBK2xxotZ
XlObIYS5Rg7+lmvbrjJgNYIK5FLN4l9fpce8jkrsSD0hjEIXF5gLKv5v37idXSBDy4oBec9+DiYk
nUNsUEBewPsTVVjXUGhndVlMrPerYt7yzrQY3+PaB1aOMz+16XB8S2aP4l8hqD7s3f2aKp9rteYl
Cu+bWEqFNlxLDwOmcTS2NBeLfQCW5L/d+Vm6IA/7fJzXOMHIzLjwipgWu9VFUTLqTYUKTOBXjNgi
Z0U9d2ZjSRIN8K0bxvCYMwmjqKLRVHY64u08I7aYaU8f7SENU3XizvgqHKzqRSktcQbPwcIeF51Z
8e9Cuu8wMf4Z654L4cpECsY3oDRLc1pfEx8Pb4KfuDId6rnSp0s6M6FhLc18BDpfPevtSuzZ0TOY
DWh42TRRkM6mQ2bOf62iXtw0cbt8DAME1rd7X+/O92gPwJtZWjIowT+1A+KJuUF7IraGJVQRbpee
zP9xc1N+Ox734FN6fZ+e6f2MdEExXqiAUaisnvQE0JXXS+TjdqKioOYN9fLwXjjvndPmM5KCLw66
eJsI75QTm8pEDhQ/fse+UmEklYCqhEz0NjbWwkV/0tg0QdkhO0Vb0Lrrzyoie4bHKIHFkH4Uksdi
hkQR/bKZL/c8oMGts3AapkoQhBVhyb8mCwgs2rjo6TtVe9gUooVAcxSQQP3W8x9z3H5ZzoJAsSkh
TV/yWLhCkhmpmfSXUh3K+ajggX5cZJh4HUyVFtIK/iQGcNLzE8hqaco6fMp/Fvh/vXtpExJlraM+
qjak3G0JNZWDzghO+m0SCiMS3X6E8BrIEK4i3GjeFi9KBujXtUz1Vg8RsdmKgk7EBa6/Jj86RqHz
8skESX5uv3pmFOqlJJ9B3cTA3siwzIW5Taj2mLKNanRlRpZlOvq6/nTtMzTH0mYV/IgmpgKoIM6i
z8NtDw/jq54N7qZnjV8deqdq/jCvlA9vkshXEr1nyW3qfiRPzwUEHE/zZ4qxai4Xwc/4LesBz69I
KIxcXFNra6aMtbELEbnaQz3KwtJP0NytE49l/oEwWvQdMV2aIkubn9oIGG1If/PXxmkDWdhdhjKc
2UsTCHALjSaK1IqRq1kkcV3aE8vMSsIXwrZP2XbZ2pM39AeT8NlbqN36sUqklNvXktVPYLjnDwrZ
IGV2uj/gsMtS94ofNG3BmZGPPm6bLzKa5tLQ7lwSVDqv/fgNDbGMnHaMp7WjMooyfjJ2gPtSTHxU
Lre/CxOCYdM0rdMVsg3eN8sKw8maz9DoE/FnlmnnUbwtexSEZwUOq+BwClKmt1JNETeI1Hn9cNUs
XZeUEzd24TeoeVf81nSFxvaNdtPmxNKwKzTrgyJ+dSTTXOrhlQh7o/duVfZXLVuUxms/mS1WMCO0
23CzPjfj9VBBillpZbvkHKZ/JqzIFD6FMvQp+UQcdSC4oU0yc3p7t0QH0xnPc0Ef5Wgi9ebb/u8p
V7KtvYyDOnlAJnlNseoSW03vW2SBAj6ncwNcgtov4e1uJmad+l+x+g4wwGqdt9NuibSN02nZ8wZG
zvrBCzJvjdI+nVA2rnf5OhwC0dFKMLyH0K0kgs/N7ZJyAKSHMZuMerku3sE22NQrHjEFvnOobqzm
ELpD6gU+DF9/Z6+pbg6/qog9kLPtNG7x1eEnKQAzIuxVF5QwB5FFcWD9t9Rog1sjQRQ1PJ/24Wup
mNm1dDs5xTChrKp1t+y/vDWBU2mC/HXXTCPPnh1yAkql6UT4FHnjM25dSIFmE/E6ZddF3J5cOQhj
J10So/s4e2N1tKsrcpyO5TlZINQwu5LoFJpf4QneORdxqrNIG/QAOWHioQCW1OkkrnldBl0bqd4B
4krV9gpJIvXo4I6pJYoZoMItVDumi32B9WMZKScycAr82Jvw010Cnji2GBuiliYNYpmXT9d5naKQ
uOF+ke9hhF8wxaOkPjCpoucLxkcmpZ2w+F6Ck+tEspE5ic63TyDoqhHtT9bbSigr7EEKKSsRtjjj
GucC6XP+ncAirmjK3rOF3VuW5WyCZsf7wSz3lwCvMVRO28Vsjl1I8isTmt3hsIjUMOfAdGnt9E0i
Za2OeOugMxWGSZXz2r67bPWEOtUWI/rEPnXHaeS3Yew8UfPCisPapkoPOpDxcHRrn/6X1vSIzY/J
gjSw/tfgGmDWa1PD5Aa0Pjo/Sh+zZ7HJDFe2YSaN+1pkZ+CU5oK4+nl0rXDsXYFW4oHP5AaTQdT1
KDd8yCL/rlOeWF1Wrbtum+LsIgtLFcYzKKnKZP/uC7YTAstOf0P+S1I9AyYJTiMfJ74YD9+5j6US
5KM/WhsYytGygBaejNY+x99ftzXR+RuYuPTMamle7gg5VG3PEdRnOKtQg1AuK/h4QUYA5UDhPVuH
LbHqgK5wCSbC5Yf5rhjv/o7yNWJ5dSOTYMOnW6u8RdPd2YBeFc1a7sFUQpmH3hZxt1xx8K2ghmUq
zYEE7VFQgyfrbTG7T/cikeIdxSfbLyjHI7Wdpg8ZirIb/6FCGxWXz8mXTmlIVK50AWF0NcXkTpEJ
Z2TgQ+lC7KSom2owd0wZKr5boU/Eu8a82Wh0nwNBji4q5H9oEDINsymqmIik1qDboJ0eeagTfe25
X2Io74w7ylT2AYoryUfIElryHuTIdkvHdNoHGpPpCydFuLRDGsHKnLQzewIrbX5En4ZPGulPLEwy
JXnHkBp9Ob1MruRClp0lVkVzeZTtGNanRMVMXnX/O1FyqRLsYmXAPqkgLhAFiqiDy5s3FJgREkw6
9bZBy7Pdh8TmeOlOmQZZV+UoI0ViK4VMTZ2k+1rU5fGF4eobL2uILf3zp6OO05Yjmp5iQnpwMXnZ
6zDW4zwK1RWIqiObtZlz9Q70JGn2icFd2JGDUAcoKTK+LsdF6lR7SNSFOjWy0xFo+EU7J+ITavh8
4WGMXqxX0KBGJCH5utdtSLcKEKTNUhItD3cbjZqfzhaIHFuayKfPFH3/w6LnYN95D2OXpFoyiTHM
IHgSGgfdlZx3evhGvpCeOT1CRQ0lHH77+as+0ekiRNf/dPp6DvlleMuhhz34/YW47qwix9y//KBe
ldwPbvP1HsmxyT8fSlEfgMx9J5U5InNzhcdTGVR8We4wCqU19xJy5qF+FIHneOFvXMlWvRaqdtv5
EiEp/rgAUQSs+1oVflWruM87iH7OodK70OAVFfel8bhHW09xH29vLe/JAxtNUTYRlN6PzyPEeQGk
o3BKzxvtPUN5vAc1zcgyMib1ZAkTA0QvQVRMpaCq37tUgaLpDhcapYx74sTvvXbZ7QHDhYNYsluA
CMmRodaiOu2/H6RuuQouqRjYZlHJu/Y7gWCnRNLVgk8MW19+BROR5dwqqo2bS25Y3ROGCC1GyKPu
d+EH94zieZum9lCN8+YN08wb50+IW+V05ND1MTYzGWgPmWzIGXw6n2ajhFexxrZ/SfvarNq1LZdL
pWj3KiroF1fdyNPYi1u9pwwggY3NwENDLR8IqgA2duwvAzTxQctpxEDJ9N19Imjwmt3eXhkrxNbg
297fxwwB+F12dHXLuXY37fZ94Z7VIXbyOGozY4vyhOhNiYRkzi75tW9dstol2GQul3VYc733tTjU
p+fjKZPfOhfBnMo+TrR90x7J7mS1CR3OUL7bC5nHRKl/HvFy1AEcQSiDslcWK+axUCiaI2piLygf
vJ0SoFgKKbK0tWGst9fCATR8eQcFEGxyJ11ZVkhbMkVkoU0TgXjVBIrawI75+N31NVRcw9S53Pow
NNFLCt984Dt+Ma6svTvYzerSkz18KZP9woZR+FZ6cIiX5xjCGrP6H9tLrMR/Rz0hAcSzc8BZovAs
EzJGO+S7YpFCuDuMoQ+K+rxMo9Inx69bi+tEV2A9+CxjU0Ofe479OjUf9KoqBe8jsPz68g7ofs6/
uPcoRfAprPJNBN1991UORu1KudAA0JxBSo1iQy5AaNz9Y1ybJqLEJT+9huF8UVdIOXAyW2HsttTR
wIANf1Aa/6aZjGDAvDX2iCfn90XBAkYTd/Gxbw2MKFdfMF8o/HDzvYnUEKM9XhyIwAl5eTErnG/J
WRHzl9bdPjRHdGMsclnC+P+Mi75m1AGY/hXRxN4wW8t1yP1np6wdzeRPjgOhFNJax2l6g0iQ69g5
Mrapdw7dC8XehUM7avzfljBpXEcAi9wBx7eEGO+dOl6hkbeuzZryg5XEkQcf+8XQq8m/zqeASf/W
ck9TENFIkezJU1O1JmvEe5LW9/cmlPM2t1a6NAtr4atPrttjAZe50Aeu+5Dzn6M7jZLcZ3lvLToA
dUzvS1Nm2iVeZoFk/kwuPSUXbuQNAkdA5NnLNdc1MIFATGEUMzaesBQJZhI/jYUZQYBCmpUGLwU0
vI+mcmsy1Jra868/zJYEsClMPF3F9yt9Iju1dgeWXx1P9BezfkfWDDFm1YFcXmbbkzPCKYgtg0Iq
6FAcBqr7gl4cYsnEX2RLQabSIi2Q+oLFkWyLuUa6AHuInk/ySsnlK7N4o28fU25LjLJT6QQb0Fh3
FVuIBS3ogxCHRUqG7OWDjc3BPQbOI1Ha5MAgEvT4rTsmWVHb1KQJKTWyghQYHUv7/OJaZ5C09Xcz
jMdA/Jb6OZPuRrekOakx34izE9wrGfineV3ZAKKo1kY1Kpx1WrLAmqxCEIOJoh3dfTNFnaC+fosG
jCxb/ilkjViHQ+NlRB1w4a3vg7NJDZth7NsaudZ8G8O/YCb9WfN4PAlBaCXqT0T1/kJ4sHnuSpPy
k3XjZ77+V5aZnI/aL7bydALLnrAmTKBANPWwRiq/F85PEASkbvGz/DbHoe7CBec9WIMl96vpIv4f
fNTI0H9C5SoppYfMyBLlCUxkXpUIcYm5xPfEgKtq5jW7i1x0G0T0fXvXnoJVyEqPusDIVtnoC0Gt
u4telVP41d+33GFrJ0/zROgg9RNsErBTHcIUgyoJ3+R56C+X5uMyUOo+ObbbY2QEuxczsoiYyGuD
JihFkZdp1bqnXyF7kKumsvtWIc/YGtbFrtj2o7gIQa1M6xGlWqflvjJIsM0TKI8CpSfzWXFLgD8H
QxD6cxM+t/qkFKQhzRBwZvsB+MXkcQtPZMPrIFQeFC5xcjpioS5TKzV1ZvsHx94Z5mqsbfBhmBGe
VC22hy/DkCQNrVszDlj7zcWn20HFMdzdGFpM0rEa6zt1RHIt3WClBh6EiVS6G6QaU6ZGmj+i/rab
mz8uZsQwmwso90qvwd8+l33ybC102eMnjVFhCLOwcy0twyA7DVgZmXCiSMR9VxxpBWJ7PGzQSVyV
BJenW4LoDZdV6fATF/1e7ovXGYUn4O/WTFAox9B7JIZUERWrXM5/RwEQ+2i04ihCGxpfRiB7OZFS
WeJMkV+zRdD4xv0rzzu3ONHbBImuX8Un5cO48YiGQacm8KqF8XPQt656OpC/ItutcuQ4BiULIZ9b
blaFd+soAwnIbwKXXTnrZNgTNcQswTBdXftPoDXaNs9L6BzkFnDm3biePDXofhB7uijIF3KYlSYD
nvriQ/csBLXW4ME/G+hH3Lyo2FPhz2BKvQuoDXiRRYT5MeD71QqdQZRmQGAfMehvcICFpYoE79st
1SAKZUFwcp9xiCE3k947HVz0MTSWP3ZJweGFHYeSsYn2nKNnNjXvjSNGrlUf3tij0vxGHJDOx6MG
j1H8ADsQs/i6pbpQeqY3k/5ybJeQeSxq/BJiZNHnmQIKrtKhYS/8AzmilGTnQOwq7jn4fKye4rBr
5f3p2kueG2aRdTt/tMRdkSurtYr3Ft/lK8t+DFby6rEJilcXDALhAfmnrzz422mUSCriyPLLoFQu
a6TC4ALBPAON15VnaleUtTjEdCnFoa2HaFFH8XZeYwjj0RQibd2IB94p7df0JPg8DP0oqtYxCAd0
e2PhWtfaieadBlXO1O+1y2vLRscQHdHprke52yIqWJodbPwFJS1OjuiiRAEA8uNRCLzOIRhHAQoV
lmCCoU4Xvfhx/XB6M6iGukhAz1uZUGpZXACUOJC8mZlDVKib54IATNAJw7aNrSHZuvWKSCbzPAM7
75JP1kznJz6dJXHdbhblt6OT4gArp9Zenbxv2xKmomMz2EdPT+Tgm1xHeza8pYTEhfqq4o98eotM
n7oKAK6oFNofpCbP54VliiPkTlMgfJ4j776uIeDhaoP69JprBGKH7v9P3CWcnD2A0GJUUIGClGKB
xHeUP7AVxdHhhNmhkgNOZ1cxW8gOKB4GC5cjlwcJIACJZZalzt1YSD/T5rkkyPGU8H5GT8gKIAmm
3EeJ7r9XkY0aIH0Cvti/3Xsj7PLStAjJwR/A2e+THiguoV4/WKzPMiYORGZdAoa7wsqKmihWablp
1RZTxvCrUndcIMf87RXgCZ7jBRHJgkw6ZlmyDNohhJNjlvglWNuw06x7Fzbs1QjiADzPwkrRuYbR
U3FpLJBRyJckMjc8zpZVSv2vZrhGtgt0Ew4xh6K+snw6NSANfFx505mZTbNADId7ilcYpSXVpdeZ
DjwujkfZx3K6/n34Zk+LhkRt4b0oXSUb2EmawwINYVTKtHM7nF2mm3RFzmUeUS5tMAytXzq7S5PD
UivPpe+z6GT7jwrUAMtDC9IPDOCv3KGBfx/REzvDSfHcjBOa1+Q0KUIt8B9rLE6K0+jfC7qSXMS7
4o7InMBjS9X0Owp671UuYZ+wh2BD4waqPFkYU4LlnbJiHvOT/kpNohl8GPdEeYhP/8OFtur91NU8
8dweQZTQ9IZljo7WKRKFlP8nHkRyzgiq8fbsLN3gU4/cpDgCMdnde9yPBKy7p0m9zCg0ZcUlP5pZ
h8d+nKK+FJ2MJENJzmCD8UIj7eDddnZNQyXdfnotqGFH3Y89txWOh4ph4pOZfVodZSLDxaVrJhrG
0Bh9yDZYAdEOokc/zTjR8M6oKwTIq619VGNCCN0HXDyelp20AilM9lBlSnZPgZ9npxzvRPonCot/
auVvqfauBCMIyBZ2bLMeMJ8CcKQHtdDmffzo7Ua1xKM36bDw6qo6N5hodbTrokVwg4vUZiuvXivo
Oa6JqVb2h8evRZytyYFs2pYWDOywV1SXrzU2eaDSuBXSnWoBWY/uPMDo6aBCvUssb/AXRNSmjR/6
WWXIFYXbSKyxZ7ZFaH8Kp+HtzmGPQzbKu8cLw6k3Aa8u5+3tuoZmKf5KONhWLTqQo824rWOrdLVK
0nSjOqO4T0lIZv87thyocd+D2M37BhcumDq4lrBozg1fDqCe0j7RLGO0CCLj8uNT3GWG8wXWJ86G
jgQDUd33JMpdcSZ265IEYV4s4okX4kDXoES6V8bLJKPMgwl+LGrjMVrr7b7r48le+mJAzsppap6y
9Pn5WW6yJQObjLS+DNLEoiClqG9TSx+WRXV2YFd7RqFWZUpNfBnObBufXvEKdNM1CXUMmgTlNdRI
W63/vExCiV4leL7zVtUbdiA2hpr8ufN6sX7tzU/Bja7JfkYsyneQQuLeaWj/KlVLVkIlZwxjKhPG
1kMtxy6FbFJ4lMeUQAmxTypO7XRlhcWtE1so2w+jbMRxXC1myO5nCHTsBm1viys1NBItuP3zNuZR
QwPzI1QAFMuNBVyostrbQaKsTEFqqKk360wpO+JUNBzgGlSOcbU6PBGJRe34sAzZh7T0b0xzhXZ/
caTtXdOzppTV/ymIjGqa+1aAFEDeSoSGsbW0tcHhvlEiHa335lHLse62YUKUgklu5q4DRolnGic2
XhQYM3vHl7Aw33b+/LrDByqfKxRYUmDi/Tg85PvY/ozZ2zp4onv2L6fza0FhoZtn8z3VSphr2WRJ
6L4QivKS9PK47huA29sHrijVvio6Tq17fMz41ohF+LfBo9eYIAfTm4ObUPYituflpoZ8FIN4quDd
a+LBWfM0q1eLQeL6yHjUDdSJ9lhVCBFLhxfHdbIt9M6OjpDlT04GJGJK5RV6VnhK1xRsdf8SrNJZ
GQ9lxyGW0BQxr4mbT/5KT8344keTDA+ZX3ECM/+LwW0zK44OYFzhMG7+FRtY3sbhrOVPs1sRbFOi
Fpn60G4IXNjfDjB0t+id7UGvk5/2hXJdn3Fc0L8vI9zzbePC+tWoaWCBqsazBbmZG1jlpPMoOOMa
g+iwDPl6tQFZaoTcy+T1RGeurYknXXRCkA1l/jZSpEakzwvu+IzAPdYTzMLlx9N5x4TPu3BVJ/GY
qiv6XU3b3mKYWxfVG6XKJXFkBwdeNep/93JXnBszxImPLw+acLS2oUAFYYKcMDhoIoEGYA+XZtJO
H9OMUxEL7DO/SK0tD77QBxQxCPSdmFvH3/AZuZvr4L5JtRKP/mqqUvAV8LtIoHjjVvEDtdFNbxfY
67hjEnySS9h2YsJ/ZzmAveYMjvTeLDsamRD/JiT8NqpG70DQfCKrLn50sPzWQryiWfu9sKJRBJX+
bt0y4ysAn5Pu9ysb6+JLoIWzB9LW2VGUqcVMA+vypxdp1IIkAq4yniHhBRunxWpOqJuA39s5fNou
OcMLOcm78FOnjWp0t66bbNDzC7kTzdXacwU1mJlROq8WiND0P4CraKl9CH5a7KHp3Z3b39Ol0FzQ
OblTQIsrvVjCLGLroTrp/4v2dL344QfbvjbvIARjtoCj7zaKsgl5pAPmfDnWAMXdDRuNVmYtKpKH
b5ceuRn2MOHBjvDFz/3tMkIS87gKVO6jbtlqihGtOVcuvuUYDdPO4rLtzN92aHJ7+4qWee7cPxwp
JdostA5RbxO4hWPild7PyJ2MVuqSKGo9bvqc90K/PePRBc/OXJgPAvCJKLsuomIYPxAG3tc2AfKV
OON7rbEL59uU6vWsI26FZq/a4vBxyjsE0ErKgNtphgQEWvSqH2gMeEPJxOfGjCLIfAg2j5hsysbQ
rfQUlPiWJyB2MprTZic6qxjO8URuMVVSPgKYU9zYVbHzM8ARhOmt8ZhSr+TZKhmu8Ub4qyVbe1xN
ciOgRF+CpTHsVucAr4fLerRfo+JzGtO6rgRF3D0cN/drVRMJLKubs7CViI+uEuycbzIl42KqCXof
qh+z8nMXGRhEF6PF/lyWrWpo/2aLzWssdTGv6G3ehM6h+sDn3FZHwIfGwhjim6zY72hbPbUqFn/f
fxTgFH00Kiu/Z7EKRL10ob7cEe34u5K2qHAx2WyR7LR7dEDwsf4lWxBIK7q/fOWKyIyG8rYgFMMg
qPJhN8fXjIW1v1QcPyqBTmEkcqPZSkSMfTWOMnINQIMhdJdPzPvTPBFPFIoi2AoKE/Bbp+rHc4Dz
DNhvtcPcUwGGxI7KJi6DxjW9cRnO7P74GlKc8ndNNNvSjMIa4JiT4S1Q12tH9eIbSzEPka8x3X9P
YRiYqFPAsc4LKbIlwUMM/PjOlExSjbj4q8knlfsFgs00hSdfeorZ1jJgdKkt1gKGkJjjnfEfEBBM
mCUc+RAsZ1EfvARVkYW2brRwTF/dc7CcGYno2MOKeR4CIRuWQA/ZbR4yTUFjauxjxZfuKf9gGaRg
XAKksqatz6st0xmy7F0VNRUDeJDUFaTRRSWrqUJp01PlSCoRj34nExahHz0Fe97HI7IsQRX5YHuz
xAPoOKbv29A1VDHwjYbvFxdGr1ixLn+CcNSusTYPGviJUW9EaeCDlqMxLaJZSueu5/0hr470hBT4
14lTd3inCYdUKHpeUDTXXZ8ckwHFfWz9v5yAoNt2nZFyw+sBLFBIgqLkBxLK4e8umHGdbY76t7Rm
9SH8G4oeHpQ0YLBrHn7QknbF/BZfGBCMXsPDtwkUceM3gvgZ0EvmGLvF54MdR+PzANrMIINd6sIz
SHnlNeeXJnPWXVfgtPWRlxUM2VmuGw4Ae4wk7pgxvsGrHsnK67c+aYXdxXmzEzmcbS3ZUIPS8Hln
IuqC7HnKusZnhAU+7sQBW7tO55V+fyMKJM9O+edtCEU3JKx4B/qoA/IG78haKgaITcjt7v0hppyc
Xg6R82nozLbyxR9NrAjRwP/il9t7a60ySKpdXHlTvsBxhKyQaBppGKhi7hphsqBws+04KzTtI46/
gFMkvI/NC81O/nU0rDwlKqNjZ0rHjz5KtXJG+5CWZDXO4orGj32YjttxFmbTLTgP24VpxSBYsMow
ke2gwKx+jq1HvbEM53Qc1duQlXVEbuzqyFVCVeETplR3L0qMqv7YSqrCL+DRiehbHfwt1BdkCvAv
CYLDpz6adDn74O15t+XfC3dbwHfB2Uyt2qkAtO7EiBIpVoeqYbXcG71VKkMpd1Ks8ZA1jcBCLYdl
ri33cPNcuDzo/DRww8uuwAQpCzBv8gew8P8ijeyQV7pnnxwb8hEGec4lgfWZKpbjHM7faLHu19xK
eWG/U0TSb5DYkePifOhr6fXBBQ2GeJAP2y4xoeoC98fRmieXitLyzLKHGaxWoPDOvaBqCu+ljR4N
KAsE9+m3kI9gkUnBasbwjR1tTdXpuItamM6kPihQjXYXK/zgJW/TjZcf9PSuB1q1EYp0vSCE56bu
XotNoQO/jUbdWK6xCFm+MEQTJ0NvzBbyolhW9wqmmj0r8VqgmBzl8upFiFG9VbNV2y0tHROKtAuc
NlvZFf2P7/OTtBrd3XzdGA4LlylNSqnpMvazupa0JplAMhw9aSJPBmacpTVO5NFEQk0FUkXGd7bi
8Xs7+Pvlxbujv7c29HYxj78e5NVLetGtsHIHNMtjRHrbxskYt3k+X8XGWptIMBWnKPhPz2CVjYgd
NB9tz99rIoGkbi2LLjqQwKbt9I5/bvgvMRxVgoiwxTBefT3DJN5DzB9wFfrG35eBFisae+S758VF
aNDO0d3+kWIsPWQKL03u+/bVcnTvz8vEUnj+PR2GvvNfaKpnxF6UFozxwGKPPw5a9gCa5TTx0j+t
CZ/h6PW9/pU8sCKtoK5jWn+/MJFXFLqxrTj+9YZyzffieOQlYhnhUvNXqZiZGE/InbvtE1Itt7os
qst3vELygnqyQyl24tM7zJCFjy28gTc6c1xsah3/bVkLCRoEgdy0SmP5LuVLabg78Jo/ukpligAz
j9axYzqsd99qeLiKEvJIdul3WkoTMrUOXqy7yyu43WTpfedqMC50iPQSTP6FwZzKkupMvvk923iQ
ZBA29ls3J/gP7k1xBPpyBFKqbUSXzALMiEtI1evdVo3bWeJrCQNbxFA/egNu6S8YlsBd7X/vcn5u
J7JNvZQ3nzbyu+DS/Dyft9rn02ujP8ZZrJ/bIkcDcX3I++YMmwcNYLeVyfZVFpfWpol6ofkoUFcO
2hPsu/DQ6Ix6Hr4DuXAZcKe+37YYdtPfUsHUxEWBcjdEDYbZHBFp4f/Dy/hmtSSE9A7FLq3YBKxn
jIC6/Q7zqNgBxuAhD2OOdvcivUnnbikKeRHk/58y1xSiG9dN8xGwQpKlg4dGBqKtcnvCDJbzK2tc
0kxVersexV75rufrLbLUhFN1WSJOl064n2nr5dkHc5DULdqHToDyZD6iQ7VgvoTpeveLo6pb1b3H
flrqSBIzs2P3fHOxR7VB367lGH8u31x6gYEPOGU8gXTtmB+tFBoC8lQOViROItZ3zgglPHzan9OE
mn3DM339dIN4jLPjqhb5kAa9nhd0CJ7Y4yDXeW31aLnzx1L5IsvPeK51nep7VViqOCO8kpMU7YJl
rYmgO+pQ+CBtwiXvddZ5S9MH2QszXdrw7/ZiuZLUPHq8NNd3nP3X8hnM88iuokeR+8fV8lxoua4l
5HPxqFTFcNewD7JOrBMJGQArbACLcF/ZKC+s8O3Y4JFuaqm54WlCx3r1uNzSDHD4jNVZquUuD21g
eZttV6JoMbSxL7yy3VB1lLu24lRmxNdQz8ZGCzkg7iUzZgaR9YBpD+4F1f8j0QlJanG8j3v34r2Y
nPEB6rIjcoYnobvDhoWIQHJzPIU5EM47TDL7XQvFkSi07e8kgqScFtgr7ekRSZuCEEBMQJO8gg4p
/PDFPI6tAk1lTM17t3tNVJ7QL5U8fWfMFIwBc5PzlyFdMxEs0a4vU3AYEqdRLCJawVCpXLYo8lqX
yyu30HUAPijjbHpc6KaDvlwlrP1Kp+l0NL+UsF9hmV80F++aYZsYiklv+2cBCuctXtK07Ea0+UXV
AN4KYNz+zmBRjMlN5MlYcLJ7a0R9q3Qz8W05sa2IizEjf1JVzSyDMLcchSe+oruZIZn2tU+wH7lI
5H/8WVtDVlJGvaGXQ5In64/zn28DJ0IDaPCnLaAwZCBpZoiYSfl3EB2FtREm65ZDUag93i+kDjLl
+eJDE4930qL7Ziy0By8wmiLjLIityFG/ZcH5yPQYGEHXEpAZonqIGWPRdDfMIlIjQ5caJS30I5AK
duTu/aMCeEE2P7j7PcDR4w1keGT4CzmIkngURRhWXVYrurjLOjn04Xy9oafixGxJ72HmZb9Ig32l
+U3043iVkfRJxemM/npGB7pXz2GW5r2c/ZXsSu8Qp4zHX5Yg7k2E1mv2wr0b6pXyLuwyEjFZ4Gw/
gOtqNelT4Sr8nvnuxIRhrpLoYMlNplR/J1VyfPND9BcI6uGBHKQ0m7Subtwh/f0hdvcK3XIXNHiD
oR1WzXcQbXvlsdfrScCIKreAF+fRYX9gFN5P+HUb4F/d/ep1iObhBZ0JEKm1ceQDB33vQJLxl+GD
aKXcAjBrWQuanrks8G+2rJjneAiedrBu//PXSlahphupTF+RdVE9v2zOLylx3OiR5GQQ//B9TTos
5bze6lvZS+m7N3b+M1y8lzZZSdxHoA95YuII4H+TFSMNEVRe6T0YAzowZ6onPPq/hCYm382YDlth
n702y5ULi/G8MW+COesUBKn0o/JI3iCEB1ncjCgV0dxq9hdHDNgmcqjajR1jcSNJVTYyw0LPhclT
uWS9ahn1yUvc5m6bV9qFkHS1ol3fL1GPKA7t2ayebSvE+pBWiF5W35dNnPMJuHxiGPWSqsvAempe
svi6MMtc5I4D7LwG22GCMW1WIIVfHWTUVAcg6hw/UBgoKc0pyRgWwi5sma1atFT+g/ETcZW7VMkK
MbynpXj6YTeBjl/G7S7/oaGt7jRm4ardH6uPyGT6TR9DuBrB+zfnMepmL74SHdAekYxdi5WIyhf4
9SE0DEQxQ2v2/pYk1Okx/5dCtrP6tOe/gFgHinl0f2Agt8MMFs+wEdMdx9BxSYWWTXdQK/XwRdEJ
LdrZlui7RKfOYJ3T6NFgnaFMEr7lMvK4HS4ckzRVI81LBFZqK/5zbZlo60Rpoiby350VZLzYeD18
h8wI2OyhZe7lWTP82c5bylrJwryas5QQzOmkDDAnlP3KwqaRRm+nzJqIAhcug/qmyyHpPHvLWeOP
xyb2b5wfQPDFwzLqZCn+OdXtCquqqZjYLSB59TDh8TSp7I64DFQBWGOuFNd2gcJaWSkZCiFf/fHq
ehkNDbHVbrABuygzA2CGAoShCpLtqHpq1sbLfg8s3uFdePaYg3dwvI268JXOx5xy/yLZt82TFQvH
3uKW97KxEeVRlqZ1P7WHeh2a9udbdwpG2zhr6JV/nC1EydkIveuM0YEK5auEV/MSC8SVp5m8lSej
eOi67Be5kcJG6rbq5X6YxkQwJV10lFOIYYlW1Gwag5IKzfO3XJ0x+PAad5FJdcqQy7pUuuYpu1GV
3TMp4BdJ4PXHQ0oQM0l7GtHcOYYiSqXVvgua0UowIitq6QL8GLGmKvHHxdkNLGRlAQHVKqYWUw/+
SAOKnCbPXKAqaN8tf4GYfBXX3254Ym/DQIZRmfVwQ/BAzUQBw3oJQIce+0XVhxSb2llpNWYF4lGf
yzAwUMFS+qSYh4l4JYjJfJBZlt4/dG3HDU4ZrpalyAbWorBl8hYdmEK+RjwHpwpOFEbCYcCE7IuJ
ZbO0gsuKXCscLGqe0Pnqt9ouB5ys3F5SDOgbi1jaHT+Y9PmhjRZ5k/CZcuc1iEHU1xuKF/EUDg9N
mwbZ6L31HgK0o5P77FbXrxzN79dXIYhz6zJJqgvTjkyL5W4DZPu+B4R2tWm/CyGSpgBc2vDiToVy
0riEVbgqtazCd+zlYj3YMQAbahITG6hByvrewqaG09jNlGd6O4aOJ5FgS9GVhNtPLLc1/wfsmWR4
j7oPYXEMRLDKSPSp1FIMLftj/5qSRQlrjDmHhzH5rq0C4ICNtvFVnMdWRT0sw3ln7HMVwuV2WMoJ
Y36RXp35DFyEEZtwu00dVU/ql16BKgphY5MobF+/y6R0y78YztKISsGXFetSr4lDtfPB80JTqCL5
Bf6XrH8QmOsgbqEnVVcfxcKVbjbY06hQUL5YYNWAzFmJ87vsMWZPJ8s8IvONzRkJ0SLCSjr6x2IK
1RzAFhcykGn+QNeTrpL6HjuItT3cgw+GVXv80knGipGCq7y8L9j6qjP7PVibwsJLmax+RyGG5GRq
91XmwuweI/oIKKyoPL6dgOh5fxje2AcsJdd2SZA18i1/Q1VPSJvGTFlDKnxL5plIBHtW2Vp1tSsi
ZZgYwjaP9QxkcxbTEGKS7BtuSLyWDHcHjr392APzPd7rgZ0vefjrAkvEMXtzdpgBfGPQdtY7H4AE
evyHIUN3+ht/FWdL8VqNuPVW3zjxmk1P2jvTR9mImLwiwMTiCyaz/DOB7LVlrYwK0YrXen+JsW2K
LRvGwfuG5qanYYM6Usv63ujeuOuPqQzIVly7yQaQP6Kd7vrb7LXy3D5I9UMuZoi+D1Q0A7Uvpvw4
fmxaiyZNMinDXP7Q/Aj2+NzwkiPRHQUR7IOZZ7jg7qhBBZ7cbOfb7zlP5RtkEXmxrVBTcURQ+dre
nO0VD1WyBwIlZHNnpJSI1GqTT259mtfzW/59m+NBYz66yYYEq5gxu0ExYrqcZK1IUKVQW5ZSPSgB
HFSZTqI+vxJWzCensSCiLFvMY2WFx8ErDujCgfEnBH8E90q+9aAdabQJm/k6HAy0HHV+EsGMvggI
w8FHNcrovA+CbnenAWH1Nkn1EXg5KdAnRYNp9uHejDWObHm1uhgUJvJ6bGeU+BpGmTRip6yACk/U
8+DbMtvJLYt0aEjUG09aS7Qo2ohzAQvfqcodCm66qdJdsKT7POR6DLDpTKv2XijtzvX99+ZASkyI
zJ69i12vQdL4K/uH9Rp6JA0NwgD20arIET/herpirWO96tRjXMWNBkBTzKvjG1tSfA1hYa7zwXke
mXoWUl+twQXaSO4qyBJk0NUniZPtMh906fh85IqIhybQOLkilHKEn8veakEMRfo0hu+m2JQwZWka
h3s5mivGouzWIeAIXDjZZ6bpTwFdCZgGMR7YVBhn1gUJ1Nr3q+DiR+gT1jc3v1HIioK3oGWSDctA
Bd42s1vVkR8OQW+DmiDj+AIeC3wxMg+cPUq4X+JOZeiugTzumzDFCuIX0HYRSCqNhqrSn7AKyyKl
EK2pL/oHU6JeO14beLcVhrI9uWyJL1ROAgDX5/FbnwfNdcNBTy/62VXXfC8n6noT9ippGktW6SUW
luNxKfyVzs9fQ9/O/tMHZtHRzJlCJWkWbX2yq6Z8N9ylyasooubq4C3yrsLKyw9kVxAanuCtSl6t
isFR3vb8Y9emh7P7dUOdceuNqmFg+cKf3uOHUTNkMpyQKxFXBHe6sjNKeXosFakAoWBqyxCyDraK
xtpFuyqlXn1bgmKSnRgdpVrDBYv2IW26eYbCu3kEH04pZMbtDHZpl1K6/sKJg/9z68zuFXgpBYvH
xd2ckLKtDgA+Xs0c8GuVNv08xXBdRGf5riCiImGvG7dZSBNiOksqPhhD6oNb0/4827TJ6EQCNXeT
86wxaeuFKj3qExYtmi/u9/R+Dzif8z/nxxGTEXjGtJnEN0/oe3q4+rqF8atY6zeZkt11vcq3SuOA
UuOR6ifQux6eL6ec+s0SPr1kBqa4oOfEcPayFlPZAxti+qdueILZl9bA3vwl/0QybBzZrvCpYFb9
69XJ4wGRYFTRQlWpaxXeexCjA8b3Y/4XwcqEm8FUBd+oN5aKvA/DWogmHr99ChYg3/St7JqSqoFX
WYvMXV1CRAEuTSI9/MHRKaeVbOWd0tLYcb2eOdstS1o8HaLWpS8y+16eJ6Y1gQAgUcAI/+9XZhQL
/92aWU9YSf9XZ+HHyQKivHukdRxCKKc93XOb39JDxqlU2FmawXJpoAOe/Cc5HpEOC367CT3Bg177
uM+mogPaDH04i5/9NzH968+P9Q5yajIm00JusvTm1TocnRUB4blwCBfg1wZzHOwT7HAeVrtYMi6s
knfPyC2qMnMbsVe4Qk/Pcfdll/cJXDJ19fl7c1+VdhkkvdYROf2FoPfXaJ56ycMsH/SwWNYUf8eh
XtJIDI3wKOk5WWCxX9NSigsmrhvxDDu1NI5tMTwFv2gWP4Dd4AozMlUiqIlU+xfEAZnzgoLsVlwZ
dtxnVqCeywu8WiyNUN5J/xcuohJMtpHgRfarCj7/Kif6nSzznpC2EBaR9ABd4JhTppso8+AZEiZP
svdBBCetChDl3yfruqRVc5zKz72Qz7L9pc878ZQibB8MV3R0nJuNb9McW2kLNXZLzllEZXw+fQAr
uRns/lSIpjebofQc1+vQTTRlDLHNrDRNw56+GLm1C55EAfnpmuiJ6olHQoKpSSctGISkK4i/eH6v
WH/oQuTXyBz4ardNAcWGGkdoKmFZTH1s+YBy7jdVZr0BJpE9fUuRw6TkmwVydEOLGtw4mo64SKtA
FIgMNhaHn3EyovpPy6D5sOFfAZwyPV/j8y+doKAtVkUtO91ZIoTqtaCrxEZFJt/gucQWtZTJfF9o
szsebW1m3PI+c5QKHX80M07W9+P4qJ/S0T4cS4LPrKZyRhnLyrKTodXv/tBFlL1Yopv06uAVAY3O
zRs2KL1H55mTm2AstCgBEJKxzjlI24K+86NM6k1qAn6f5xhmr8BZG77tTyX81ArLPIb5sjGb/Mmp
S+8LhWlPZyWKYCEB5nZKKj636ys6pT4PJiojAsfHG66zSFTV/B8YA+pZuxnXzFQIAnbzFZwHcM07
viaeb50nbHdvGt2qRd724hVDz61hJj23uFVf8IIgOniH1627E6JLMwjKCJ/4Xjs82EuKeOrD0npS
ApPVJDJfkGB7+B9Tvx+arMgy/2tniaDq6lFy1au23e1ZVzgC4UI4PJVg2gKPO0QzBwSvutYkt0CH
cLjyaHgs9z0qJ06NbjKQeXOy1RuLfNJjADm0Oj+nJttnkUe3XNtROZ8ORyEK+AleGeLWtTtyIE0S
/TOACBe3A21oqw1TgsrjsQYjL3K5Wlpy2fyk3NKLJ8u2ZlxThWkauQu2v5ovf02XrAOEESi+xYpI
n3YesOzgGop3bQLorMx3MANF0jV5dtZB2GS2z1GoBhmhw+rYVx4YoTp5MMVQFg7HPY3ifwOCNVkU
WytO+Z1ixs/nXLTbDXARNlUpNRPbcraLFgJXNdvNcheyj94hX+0BiD0dDQgPGRS+ECtPycx517J7
SNZZFKDw/hjTGmE09CHo/oouHZLBxrt5g/ZAOQde09F8ORFYCCGkcykPQ+wkljz/kG7EFIJBafhK
0nTWUUnphY17vbQvs1zCP45S8WCUQxMck7mrTt24WdKGQAM898MJZUvRk5XM5ybe84Nluaxg1y5Z
eoh2HbO3AuDJm3Z/Bmzpszp06nU4/MY2I69vORqHfucraaRIvyJxtBD8eT/0iUl11W9DhxFZrlu3
9vprPtW6jPWzAv+yusEf6Un+kCvc0rwW+SMWbQOkMMaAo0iSTkDpNobKGEo1q9H8+bPJOp0+jCgS
wnV2dq9CQFF3dXFQgPR0QeXW4s2EcZPHtNDGJcCuHeIXoS4nLAX5+rEO1GAw8w0lXBrVjF10PgST
barYOIiUjzH2xHbIy1SWWBwWLmM+nN76vi16D2cGbdxR3VanspvkH38dqflh+iLFr6VmLdTYnpav
VzMbuZWEmAz9f3HxZxJjRMINec8yAC9jO6VCVIg7DXgP/Cmi9GKnw18uopjqBCDo/Bf/0DxyN2dU
11bqYiO+LEs8CXRHwPEuaYyJX6oaN3NPgZLAHaNbEMjf0MuaKLOMXC3yFsOA2m/dyLCrYT/xQCFc
iB+bac2ESvXsTbpcdq074wHUvMzug07JhsTodY6uu+pYdeEHnFhFTgXXSCKvldLVNAo7nz7d9aGO
FOnAGeq6Bo7px60oTZGUIMUH/qkiSOrifKmfLeauO27KApu4q6hZ36vSZHBi1itzLvapxG3X2mXV
r4bPyqp6UTtB1WXIDdqg7BWnH0gK5FQxbsFQnFH0yrMaMYAadGyT3HIGX9KpsRDJiSvaaQqmQRnx
9m7l46I9T48/T3PGTnwhWGjEwAWNcAnD7L+gVH+YMOk5avgvHKkSUHOC1mOXACepXGk4pAHCxOlm
oGeMt36Q3ybCTvD5p3gPd1UpB8gU9gjKd7td1oqh78xtWCc0YFXi93fueCni9of8ATzzUsQvSXf3
95vDXjz67gyYOD2yKpK2ljD0kDEP1Uw1BUPK4eGlRgjpBcJBmtqBwZR8AkLHHa1V7dps3UxX+NCy
0Mh3MCon0PnkD3Oc7H7rNjrGAbSeLJexxhgX74HfHR0kXkClo4L1f5t+3WZ2+xWbzxqC1ZUwITIp
K3nx+r0Vj0/FLhXHn6qddntV5C5D+sjb6ribdH+q2sd7lXPloYymw9f1OJm43UzOUjcQolB/Kfaq
CSoJgsstZ4Ii6jYV4/aJgnzrBxo+BPmvahoWICJzGyXA5uVjUEmdtABlqUkMiZyshZWJG3syD2kf
vpBlNIDJ5fjU+gPrRcnjs8RZMrA2vmlpphesX/Ex1WK4b//ze2vuKUpVFJ9h2M/jStXFo++62tKP
Xm/Ew+xxZ02lxiVD4ZKbkGvBm9PfHyVv296UqY5VbvXMpI5nm4UT+kednkyKOpoQta0HL0Zt2RRx
Sk7Trb9Od+mP6qYh6RvZ71XwXNhFjDb5DAn3HRepzCqr8y1Trw7w0Kh0jnq/IxLUrSnrLWvJfudT
E8n3Ysev4lwTaJpmMWZBwZ1mDiShtvtBscwW04SEU//k+J4Zmhbopoz5RUbojhL40icWxJGjuRKL
AEZUBOtBvB0gOAoIkjcEP916xVqvaeQx5mCMWn3O+6TI5Q1wrg+tYaEcpTRgGo0A6pswM8NuDTzz
LvB8L5I9OdR4Ij/LC1H3vZmNREAywcZBH3eIFDNPCnQTVFACOoCyDhkGEruz8asp14rgcwr6DvrV
g3fLc9hPhJHQ44wYIfBSTHIPOAoCLAOEUiOV/ldlVr+1wfIov1E6JXLPtfnClDUQFiVPhM7pXqCJ
qc6F7guJ0BT84F2Myk52EZaMRfoYATTVyJD7E9auModPfWuoVUnyVk7O35FmSjrFgjWdJ/vBbJzv
c2ZREOe8/yJjxzhO2ZI9xZzckxY46qCNc0UHJZpc3ootZDXexivZ0ZTYwo+rhLbaQ0YJ9j+KBlgC
KbxJOW9Ij0RsKmh9W5WSmmwjH1veOpD/pHYU2lWwrFaOeb53oT9DVjX58WlPRijsAPpfz0BxDbIz
e/aS5WrPt4FN+WS+rsE21Xv+bWeoNIdYNBC6OnOkkDJzXiFYCxJWQhrDfZgelc+V1ciB6eK4gFaO
cgEGkKr5Ibaf67rrV3cVC6V/+otBFktKl+6b+2xAtazgcwiLig2ihAvSd3ZJYA4o8kjzf43WAMUW
ubmOqm+L5ehu6XJhK71VO1u4yKcyyZ7wj3MuPjPDYm7dgVgIMrDwnb8OaKdvPgYSn1ZniAg7k1kb
CDnkVw1BZxzgrmbUe4BE47xTG551nhoASehM+rNCMiOnWAcB95TlGkUbeamc01vdCQF0ZIfOfNrT
9Ayk2snrGUmX+iDsdTKxim1UAy7OIvEX+inHQ8okyy3hfWLu/zoF8jTluiVaqWoMng1osmP6rBtR
leGTn2PpEF3cF6V8v2uiws+y/pCa5Zm5cCRfZ6aNgFNm4WylerwZsuo7SkF/hZz2eSjZ7iAyD5fx
x/Cfzuf9tPFYi8Yb89LEc6kIFAojALNE4pzPdQ3UBfrI9MSXpKjFTPpEalRl3BmT/Pj5jcImDv7g
sR70fLuawCO+LGRm8z1lRIGpXQkX507GMNiJyCNhemTOWZkR8+m2HRXLaTDT+IzfkSCBDh0Jx1FG
l8GXHzgbJAgDrgV9AaQn4g0AXV5k8dyAtaRmANQTlH2V3L8A84+oW8RtgEIn+M6qTrl8YIC5sOGb
ar2Twcl5vyB7EjIqHCQty8Y0ahj5apRkIS/gJHIQzSZJs34gnlDVHugcIXbzee8MetHAWqoyb34J
hyarqQ0iaAo4TwHuoR6XgxK9i1FLAnK35H5PR71Y0bSZQ5lfgm5QceCgQNZM97VnKrj0QHhDWSwf
7Zk2nmEPReA2gylwbmD3xSUR5Zec+md6OnX7rcxtPprAx9j1nkDEWBoN32zP9sr6QI5kvw3dxTH3
OGnVTB6rFeJaQMX8WPrXvvMRE5+AsPUL0S7fAGgXaVhHp5PtTZy/0ucgLrUQB/e0fL+ugw7VyCcA
YtloPb3VX6FfpG+qC6h/G0Lq86Dx27P62qCqIemJLB0uSO7umur/1OLxFhl64H68Q67ll8gREaGo
VpWj1OSJC/t7m38RPodyMjP1w5LMY3lsbtqlNdVfDDsQ2tIa0rQkWLuuZRzHKVRRdYKzfB61ufrp
mBCfUC2TbqOjVXA4tFhdlhGKcHxLp9Z4rvgYenje0PpMBk4dHpC07d8AaXJgyoM3b08L/KaZamJV
xlFi2Y2nvXS7rP0qmjaSNXq0mA8BVeF+cK1K29IHllI9MaTHCe5Dav/RKVdEG6u3StVkYQ1insoJ
nbQzqRe1DDSh1jNY8eSiJcmV+24nTZJDmZWw0Cp+ohw9jdWlN+7hQ1wLmj+Ftk3bOv3HlurffsA0
QXY/cKSt29PFjrSdbR+9UjLM2/eAAYaeTS+PJg5ZhIazIg0FkkMbB7eslRZ02AYeNoNxADbCFsYT
eNmq8JgO42FNoLR42ggiIf3QI1jnFHjY0u1Y4qQB5Qs6thfd1iOMU2tKSzPtgXxjTHI2ZALokxIa
qpWoDRsnXRANHbDT0HZU4gSNCfhN68NtyFzChtW+uAKx6F9mVBDad8kXyf1G6K1f/VNWpKmmEHHO
OCXPxN984IOzaongGpNdGTfpMefTgiJ1B8ydIMGcJsiNN0xuZMJeEh9M9VXWHcs9UwpNrOD1Mjbj
g8LOl8dioTrbbqxd4ypEKI+ZGyvf6bnqeNML6zHVBAF/PRtnPxHfuIeO1rV4KGMem51TFcK7k1NK
cwjsKSlYugWmI5m8CBZ3ADtzdsTMbA4fdORv3ASe2HFajc/TOUgnYntV10RktzfAc6TvnUKoTm75
qPNJrcmVI7NJBleMfVl4NqoHbtCXDf7K2bZTb47xMQFIFzYTonp+P62dzKrH7UTblk9dmoW64DqP
/8EzAAPNBIZjD+0fZaBYKRimJFAYrycIXcmbYci/Op9Irk7XGtlIrsJ61ZkGxyu/xAk++SOh79Gm
d0OOrHTXzlAiods2mF6baTCJnzZrb17+xNfDSqnLUJ6HJ4o3Y2DukBWmLXVBHwleYMVS8h9l4xUM
NyGqkVV5kh01CIwmdx7pvb1ebJqzNMjAIOevJRQ9ht3uYdGVzXJwmGa85UQ+gob/X5/VWrctf4L4
TMpOwVFwIp3yYanvB+8/aRN+vt8IM9dXSJxbPHOkL1yvNyuuQpmP/y/RYrl24m2V10v1qp1F98nD
PltbM1EDruir+WHhnQOdgqYcnpSqRFq/+f6ELyyEliKLGbRz4t1ofz+n8YIpZcCq4PU8e1iJkHbn
H8INJqI6kyGL35j9+HSIK/hKB1p1C8UEQVuxjdxABJa5VoROkUVI8WBvMJFCWCP8Mo4Syl0joARN
vjopJYA1Gp58GTSwZRaVAFXaztLorLHBKbpySQcQSwdw0uuH62LXWYGs9gDGc7rsZlape4+IeGM4
u1YQWB2lr/AiQDsgY4cpRZ/6Drj+p2s0yw4LAxAdN2YWfGkYHfk1AqS5ghgDnI4xyY8RX1bCjdTv
tfIqiFFYRcr90pHQIEzgCrKQu709Q7QBXojavQe92MzOkePdaMkb9yD6CjUmBHe8dCVN9jst/8Z1
ZPK+MGS8lS0NCS4x3oaDH67RlSS7gvY2mE+5SXWt3JFd1hD1JctG1LKItKFkBtMFpnfEc5CxgyMs
Co5GLcKA8Mf9gsE03tdpHDzNgYjgxaoKk9HXa4nyg6chNzlMohZay7XoIdlC2aOc6DcWLHhQPxg0
mZIZxukLCVFzsD0JED8MaMR21czWDUUNnKj5EH30lUupNgC+h8YvSrHdeOIswcv40EHVOaXDv7v7
mxRyBHWvCBIIZtk4kAXgEe15aj61spCsxXjIefVlPH+Bscz9X7XU17mUauIkjG9+pUX2cDBsb+r1
ztiPf8WLkMyECKAdRu8NjhGTBBBh5s4g0FwActhu1Aw5TmqjxgTh+Txv+DuUz67+oqso2FMcF9J+
IXNLekDPVsHGf2HH6RvJEeU4fu4WIr1WWUom3NZCtolHpFj9E5TyQRVa1HKwGHekHrQPBSltLf4J
gFJ/IshUT4NDvlqmjWoZUjE3a0OVuEm+q0tMVAjZrrbDxO9fGBXBQ/GDtWVtkqz62vxgvC/anEw8
1QLUfwLP1AB13Yk7xekS4GeTE9Pna2jMr4Q3ERCYAt3JoDo+jB7wgByv8u4Mrp7CRKrUTheZdaeU
eHXlu+sGY9+hfj51s3BUMduNgfYqzdRixMExWdJ9liAxdVTagdSRgLW1dKRw7SowQQV17OtKyg72
f3f9vZj1g+97x4KT8rJYuzx0uQdjObvDlbJfNDpt7bv/T7H929y+A5nU8ESHlnc3LSX8P4Bsx3Vn
pVhBGQRl3+ZIv92KTXKGLkIR4Lis8OHL53kLM2bHoRMCxy2FqP8Gz0VgYKZtQeFo5yBC57vUoGMf
cBI3wB1xgquKDm/s7UXwHxjfzV5fKXsjQcuFVA5GuFAtn0JuFXQPkBvP8bIN9NmJdcuYIx5QXJ/K
yNzGEAUzfG8JDuZuv6Rarrc5iZiGuJGqHfkdPg4BcnSXnrz7ZKWGzOUn6ncnqT81WvQa5DDlD2GB
5fBT/HWl+3FhjxhWA0AFjoEKIyqFFms+CSZ6WQivPLfKGosrFCEj6+TkFx3ogaE95FJloLLSgt0Y
8A87hOTvE27wdKWbZjQwh14r4wJeQFeFrLdVnsZKQuD5Hn/+Imld7CLU6jMBHCfaYLT2oQRCRBQV
s0Kgu4cOcyILd2Tu6q9XaIw0hGoh5U1cacubNog3P910kkmWmM0l2dy1J2LMPHTsKhCVPgnIQFlo
18uIB9mSBmSXg+RPM8zvXNMiVcutikGXumKiklDcAc4mpp900Tx5YGHaPupfiB/LaQKz/1PskUIY
1Mp+AZreWCobQo7Ot6Dx+RGxCADP1LXZ+MO9muichl/pymaqW9Oo95TWCTUZJAuX/PpukygQuoCE
Tq7GM26Sd47ahOCAE+q3FOvaYbqNkZ2EiAPUeS40BnV0I53F+SV+FYZDlLBAqwnYrKSAqpz4arh3
Rm0CFSkFiRqxaypRBRof9Zs2jRdEyOd96OwDyB2MEJ1QYpUdyo9+f8kuUOSP6WOgK568trxT7DoC
fJtK+5TDSG1bmr9rWU9vggrYmjXeF4ojvsfabUdwAPbeWmh+7g42t7ippSMO3xaWV0dk+84/tse3
aXIgMCJ1H5mVFich1WOgVhGMlpeOZCOsF7CAjqTvbbhXSvekrHcUnlfudg39bdfgQtlJBjPwDpL9
uiAAqbd8+vRd1JXabl8JqrIwDeUvRNuOOx5aqR9TfwKrXa68zhgN5g4ShFjoFn22Snw/CszpdLfJ
BXfGzCoIwCc5ZmxoIH/MBU/Zb2RV0fDMt+IAKeLBG8GOGLzsfrF9CDasFKUpUQLOhE0L5KEJL0zg
merT8Fpy7sQqMAhQcVD8UmKovrWmjVI34MfIHluvQI/B5yuG312JmMTGEKny4b6Jn4EuOAfNiNWL
/yBrki6qLw95ieEN/P+7kWSv6eEN9vd2n09KH3jz3UDnGkBYRDYGwpNUWlsUsmDc8qCdGszsPGXm
3QmUz+zZl01x2v2qG3X8WNgtvtSTQ2raYKj+sAkqRMNr0BPSdeZHB1+SBVWRMKmD0vba3R6kpHBf
euceB28jYQOv87KXLMIeI1K+NNjfCK2R33kKkEfhKNy6AGbVOMBOaDCxx4iifkIpoWqDBIGX957I
sWhF1xxKGpvjZHC4YQ8zZQDetATVyMKfQ5Y/lA6TtOlIcdfFJN70Mzea7JwDHalHuDRYWJ0UPAqb
rWeZnX/poHH3acAk9FDgWuJOCJ7Gl0LzNEPurwVx1d6+oEdW0FwkS0hEKa3YFLK42pybNpAHhGAw
dvS7nu0eznpeVo+f8vWAv7GPxIxw8D5MQ28Eu7EYYDMVACU+rC56qJidxNsi4EZgsK1DRW5gSZoX
YFXWZKYWmT70QyQtBJpf32SUar27HMLaVxd0RHU3vvjXW6brPJU+w03TBZsuH8B20Lm8aIpYm4UG
ZMQ/cWBTVVr5/zU1bghdPPTiuZY3UVrnzoi1e9JHnBvnJAsigCpywmN4KZgQnBSRIojihE1txwMM
6fnM2E6P9y9y1vc58TmbgioQnnh9crFfI1xJw7YOz+HzaMQgkVkKEvjvteR6c+fENOMC8drLQu1J
RDFFlQdpSpduO/0YsPR8IG6h1PLA0xRfFL7LnHndwuvoL/jYeW9h3GA8l6XT4L5cAqlOHqLq9SwH
kOcs6wfIiJvUpYmh7Z4v+e9VQoEOYj08QWOlJQ5Mwpi/Q3OKS2BTq+8vy9rfaxpMbnn1ewjSRw7v
/sWZFn+1x1TgkC5J0sw26M/Jn+kWZo899pFXmCvhqJ9O8iYHVdJYks0A+KRy7EvtXfJilWPeZ8SK
ZyWQtMwi5wnkto+m/9DVz1d2GPd0qbDDOhGhR07jY/BmGx8CEG8xrkiciSOMQnix/crHHXuMBnSW
KQ7qAPrzmD/+p3Pm8A/uSXaI08J7R5OILHTiUvn8gU+Jjt09GJgo5B2srrR62PN0pRXl+yr4uqca
IRGlWYElEiMzZfTaZCID8MJWJtnjbNqwcEXx+IZ8QEtSbygwj6TmsP/NG8jokqNc8mNEbj5Y0NtZ
eUe7ELuc+q1eNbQM94V9Yg3wjTeQ+SuRQafE0dRg0YUtvfJH4mmAQi3HMCN95t9f1LXPZPTyTf+l
RzwiQfWlMiAE5A+2SJ/bY4+nzXIOQZy+vHsL2JnQ4Xh4adkLWO6uN2cuC3k9/z++ULvScGlDlMnF
6VkRohc+4BUWaSIqgsESUmGEtG6x/Juw7EkYQVhajS+RZ1b3qZJeXGfza1ayJ2Xjwl+iMGNp5Dul
IZBUZ6mbUn2rHioA/Ja+NMpaWmbm7gIqmMCs4HvGM6525gWnUV2JjadwoObR3kwfMOzRLjd0zqIq
JQl+Jr0hcPeT6OwftiXPT0UPSeyL12DM5VMG4ehuUyNd9t3Ms59ppV90K+CvgvmJcvNWqvdGy0Qd
4pdN/4QEAeCntSjiJgM9Yy0itLzbSlByvO5559jjVXrAwSSPsTXzrxcvnlmDwgp0GzNkh92WLsI7
ss/xTV/vh3bIBmzZjJbfyf6etF2P4LBJESATrTkZcXaYUx8FpdT2DfFb06xCbz8cGjU6DPIEAKvz
2svGqhkowQKYIoAoMNDQMX2Vp3hpNF4Av0nAMRsX+mep5Q1Sc5bT4lKjjR86t48eWh6qNl79L+4C
Di7Bbv3vGv37llnmAlTnjVVYJArN2Rz1U5YmIs7h9fj1bqN6i2docSjx91/nRsdsLQCrBShGGRLU
Z3dcjmpw6h4MnIRtP4BxLGrzr3wXZjcZV0MYQ17LnZasuzTx461AFDoHTb7PGjq/ppaks0KyeIUT
qTFVBV6owZrGvthjvU3ZGR/bpwI4P/YQ0nU3P5bvLft9JvbjbARQdVthN2o7sqYZ8olNlwNYpZ+g
KV6j7EzQ2b1K9uvzydXMl++j1BnNRki+n+Kl9BQvST7VXLLmBDc5x128e/pm40CuuG/CWId0cMdx
94I8pkUzr1Jdn+18lWTAoaMlS4eAst2cEzoRdYJMNrtVcA6BT2jKEG9HTrBr3kEHg7ngcuLTFqFA
peDeNPfr473jXwHQ/hCE95KFzpzF7bNWrUK9cJH8TZzvcSaCQVtho/FuU3qqUFRoV1hZ50fatIOd
adYaZ6X8JUNnDOd7+D8pa+iY/GbgQpA5yhD/3c9fzyA1547amG/wPVbajKeBXUiYhWk7fcZWMJGw
rgU98qVpf+cIBYz0bv9lE1u4aI4NTp3ZJbl6U27K2N4ARhVeQdoGVzDMSlbm+DG+OQMeovs7a91j
oYZuvPA70CM6EJUKS+vfE80qk/inMmbL/fRm0uER5bFdJi9AQ969C6Gj04iMaCj5xv/7xqq+iKqt
yppPAnM65SO6lD7YAck8HREkWNFNEYH5FND9xI02zb4/TpNCIdYfiEH8wVvHjMHfRUlRE0CbgvYR
pM1yLc9jGXWgil5LYLcPHJXkxmsFxKH3TUgD/VHNwGr6SXakyH1e664I2ZMVkBd4ZtQN9Y3fPB1b
cZbFxsWvcbQhYTPRw/huwmS8g9t3JHO3XSpsg0nJO7f2f1oIjcdMHEQTNVxnLteoP8GA6DsfSSWZ
86czX1MayQevMB/WAwmbDPI/48TQUXzfY9KgXlwJIrtT9ofpAAJt5azPTaB/YNaQ0CBEDfvuzWfr
eKmv1Zwyw5HN9aXuyh+oFgNe9fZKpNlbxNyesURtaNygC+qxOex4iQ+B/t8oCZFPUbXIqVj6ey5C
h3gx9jU3Gsl3nDEYaserQF+fwXxGKCHADKI9KMDB1/Ye2ezJa1VKkJ5s0HCiJ6gHE50AtHOxPJmP
l9UpqE+yv45mP572kDzCLySp7AQVxnZkIzLcZ02DdDAUG/6l5AkEBd7gutnDQQga+X0cb634BDNY
haKFXgiBJUZgZuhuVeN81pfsjQEVhDxTLylMVDkhfkImcEnesLUOT5TOcISBDEcVJeq3iBcA4/o0
svQvrfnxffQaWbkqLHR1pV5OBSQVPq3uapbp2c0o13+23AQz2JMCOOuGlvLCnUDD1zZsT8HVZkfj
uxEAB36GJfc5/Rj+Yoo6jjUt1KZu9XQ3dqo6nc+AHMUvzIceiHXADzFbPCsy1Uf4p2/FceIkQjIY
1daQWiF6+O0I1U0aKon2V7wH4zPOtw4Io/Wpra2GrJQzC0ZCwgoS8bnbwrWDvu12b+HDrJFpzxIR
BJGhNhsuUewcXzPY7tW1UyrpT+gkkqnwiMWhTWNNKr4JNRjIcJ53OwEkSREyCNVJP4ndIzVFeaFO
ApCNB870h8rmc7rU0NINXH3l5x94xn9jW9DyPZ+dcFofDjnSFhFR9tinTIM0M2wY8HSJGL5zsJDR
Yjf92vovCjxKoKep/yrvyLgiMoWa+zn0+2Ohs5bHDgwEKASQj2IJq1vTHUN73A8FAb/vOiFigX7X
fZpGijF1Ejae5TbRk+LIOgIjJ8nwjVnQEmdS7VKE7w/29SudC/pfVACn/zGjhNf/6WJbeN8vOz1M
Rm+GOO3rcHn9Vr7rT+FjYCWId3tN7KeJ340KCz3pkuOqUiTHCiv5JAYPjLMnizClZauQyrj0Vbs6
Pef+zhuwWn6p3iM4CT5yowDvkL6Wv24mnC//VMbb2jBFr3Qs9MldE368nksWDqzpjnRgBw3nh7Qk
8iYwhbqpxJ7viJabnP/w/IfhQgti+I6kvf+3iRrbE7JfpNXyEvCzP7Sg/F/3Tg55zKSqiIGieeH8
bNolq1r9xyDqg6RqcciauBMYP5Vt8St6khlopxMoHAu7yXXYFjNddHfupiFqIWpUrqFYsFZ6+huN
7buyfFg6uZMFW0KD3Su/UYjrknBrWQp4qbnT4DPoOXdF2NEQrY2MljDQ2imnO7uV1Kqbebd6dV0Q
wPnC2BXiIQyV4FgSeA5qM6AwHZiDRScWMp/Y9BWirHpoKBXrkQXhwpiWVnfRG9dWNpg0YLpQfLKc
xVCJGURUwrbfE0BYAo873m5Pq2k1fk9X5CEVNEr9jfwINSZ8F3QeEoe93DHTaxduKg0K7bW/YZLJ
nPgPUN38eQNnN4CNUCmv66A1mAY0EHogFtkA7cpFQtOqK8286Ww8lCR2AT38llsd47c96NjntM7v
KQCcT3Cbk+IitUKPZ+P17Tv4o98GggovGVepIfWurmlr8ROusWW0k6QXbMaUOHxNwqTOfr+tArV6
SH3Yc6LFcutbdKmiLWskvhQca/i/yL4FHEg+Jgw1kQFAaM81o1ey0YP/fu04vZSQgyjMhTxm8EFL
czeRx1sZWbvkqiX7++Ly/Vhx8HM8Y0oino51E0US0mLrOs7tnJJsFdFRwXRAseBdv1DQ7TuHlMi5
wvgZFrpwZikGWSpeTZ+ddpAFl5vb00YhQZGITDMfbCgAw/onvzz242TfnPi7NJ3Rx92ZVSRgKJLF
d0s8yoy8vhK4qpoVkW8kd/PSDBz7D3FNKiivT7Qk2n5z257WXwQFeLphtyfAET3aBKJ5y/KRKrKz
UqIU0HnmKdrA1NFwn0ooQLjFyc4QnrTWVQ6M/Mgi55KRqto2QJYeSVJJzlKhmvjwZp2DEemP4ho2
Ybw5pb5iAF1F0zYClsYOj1tisSMDSx+mTHB3wf6KvbQvN4lXAiME3e9kviID2OfDuHwOTcq71T3n
cCa8R6euxuYNfEZn1ONmuYfiBo6TTQvmmQCoZTneHQjb1lOBmawdUK0E4OpYewtB2s7sfuiYMAsb
Ce5K1v8l8DVkSUiAst1TCmq0j/6hJfT4KiGMO3avMeG+aHXQAYFUKw14fAt2iWxMcaENy3aprWXk
MOjy+SuMvy0ukGAunBIx4Bb7rBIXTYO7OKTkoQ0FSLjniSc4+t6wkdTkz28NUchimzcPYf5HG01M
c2fCcBV/Gsj0v5nwX3ILv6lPpFxCeAHPypJi6tznXQ/3N2bpmBlWYX11VUdzu0h9zZ3wxOQQPExa
+EoTcAxODjTcsXWppJ6viXN/zxlZl90WP4JwN+Xy/oqZS3eh+FLSE7SQ3vaezDObpCKAzkyQydtq
CnQks2lKn04Fgo2r6W/NvtvTr+mYEwIvkSK/K6FQb2eCBPOATD8wD/M4EjC58Z4q3Lh/wNKEVgGe
OZK84iAr7+ig6MOLYe1lM3SjOGID+0XBjE70l2OqKYwmXRtIosVr6iwqz3LOXM7LMvTcKdW4I+FG
HI2b6PoF6OlGLJrvhQNe+6GTu9ILoYaY5IIMAonwcMc1Iu3Y2VGUBMYxY0iZkky8Q/u32+5DJmQd
0pP5gxNN0hUpiKhHunXXADptveTn6UNXlWP+UK8b5foeA1WerL3KdWfhCQTP56TRkR1QMrDIvxLt
1wdL4+UBixMThyxWyJglIoHkLzNAjyZMDhEdzfQxosOgm6J7QEDww6DfEYJCiThf5JHYcYIO2l/u
zFkwGS2TH7N6GYUjYjBCXGdwMOsN9JEOZM41mZG/idkLMXXvFpAGj9xP/l03tU2lzlKxS0MOBv9e
gG1wwVbhonBKXgQWDXZZF9BXItscj3VxR3bJA+JwK7Eodf5apYfWOcQi6ZwJqyU6W5DwWKKCIjY7
G2XsFUonqxtraJzPXV+jO1SZWB55JbytPnux8RM39a6jRvN5gEWWfCDC3uTsCKLxj98diae2DI7y
Ano5YcPEzXJNgibrkUxOvD76CZHOVe8GNwC6SDKu7TB2DqTwsznXrs+Q7SASu5NXdphJrd368tQb
69fksJON4T/cbdEQJqze6OEzJDMR6GqrNoLGZ1u78buVlgr0ZnlN4CjcyMSWymm1GC2zeTcfhI0K
ZkzA1kCPn/sR9rerTtCUCLOqmR56FexzAHcKu9+yI8oP59O5XKhGSj6O+a1Wj8Dunvht2QB7+B6w
aSFpKThvz1e1wDLw9WJ2o7XVQ3yocS80jIo8AF64jPd6mOrtBaIxPHzaKFCuosaufNEcq1JbngIH
dDJt6QveVxOgJTASgtPY9c4fC4B/iRbnUdnLERoq1dRWKWEWnBTXashtiDmq29X1Po+ZLfqc69dR
J4TxBccT18/HqZ2YOSOJ9sjrHhojCsHJsKxk+Q10Pa4+J/fpvYBqzjpg14I/Nrg7+cErzOSZ9SGx
NwpL0lNab0PuQDqT93nx4m2jvQP1podrvEksLp6gGL+kiLMKFGm8CqfYfudK1SfFpLOpOksJab9T
ZuE/y/BHEZbtmFnotZXkG298u5C+GugXWOZcuK7FGvXYc+OC8HU73m52ApK2tfMUJox1dBMD8RYo
CE/0zeD27rWImCz87Y4i1EbKOGa6xhayappgrcsqdWaZ+X/TZO3lBCusfd9Wkdjwn3ZQzUdmzLGc
cp24oBihPoofJ+686utAi4rK9fkpiT6RXGNafDm1aeAuwwYyR6Ct84IUhB6oDrNcvkFeZ6tqtXqL
JnnpEpj8Qoh6fXY5dQpn1JAx/9tyYAM6CWfeFPy21BwnHHEOPubf0/HqNLEpc9qpkPQN1w5UFl0K
e75FrcC9XHK97LrhX3xgiks+ERRgrGP9eQZ1eZJMSV23JgA0FPROWPB3epS3Cpt3zJx5evYYg60+
DNQx2mln8eoOO0AHdLWvRMXaNuCfdh6v01GPFPNw+hcP8AApUlA05fzuUV9O6l6aEoy3xcZSi29T
XHhXArOhGsirx2s7copcVBX6Y8Gp3leTdlKqrA4SSbkbvj7EXUK06G14pRg426mL03uFjMK8btdQ
7LZuRbdCmbFW9NcCY8ki4v6b9TGBvcW3MoRYx0fW/r6dblZ//oDM8ivdkUSDogIoliDfAn18E9Jw
EM23U3Uu4eSKkX45UeYpKkOHA1iGxi6eXE3c7myEOpNgB9aD1zUABMaqPbR+3JDoie/yT2pIoyHf
I47+cNwZ4fGYzzhGgmzDrTc+xr644lTsEojO3bP4Csb6jGFAYL1NVNL+WPyhy0Jw5i8/dOkj39SH
7pZcBU+CWZoebrLryKSXpZzrgsQThD5mmIn7b3UsDxzrQbCs4ICKEo6G/UXbXJ5v3Nk95DSf4ffA
3wjaMrHwXBkKkmzx8/4Vk46SrRFXeNZAdzLh9lPwCUimPuFmX8dJNkKhFD5n9pcvCXwmfxvCYh8Y
2QsMQKYGByuEeBECqz2sziga0CUmo/6uV0GrTbEpyXNZIP4yHW+AOAUOY10Gn+aVeeiZYBJVkV7V
Ph74+tfPYp3FetZw77Dr6AXo2Yozx/WeIpdB1l1KnFXbmNghkVfPKusRct1utmyi8QLub/Vo3eBf
H98HM4BNQaanKp4HSQWgE+5zCeXZS8b0an2hTCmVELmdblOrgokIPoKzZ84DCngMOCLtnVexH3xE
qOboEhrB1sBGB5xWyz/cUyjehQR+LQc22FW+NOkyxLbkoW4M3Yh2ExENodPtqCKUqobKSLLOAjD9
tSJAy3k4hm0XV1DgQQHHnRYwOOZPP1ZXU4K/3hv5fxuvN/dpXN9PmMSEhLgWdrZwGJNwHSJ2Mvxh
5tFzlYEFdqjUBp67tD9uk3MGfv7HzADZnj3EkVN5OalgQs25LaCFhBHElB1eifoUph7KVB6ULf6D
MwPLh1JM3Fh096/sZwHkNwROiy4flAE2LCb+xAe+WkOmM0+40Hm6SkCWfNXLGuHYieUr2B2YLnsM
+VwHdWgiQHbt1VO3t8/4X01X04vgUKCM+muPqVhk8Ox4Nr8MY8Xvipnp3aiKrCV2+vnqJp0tLKmZ
oq4kmJyOjo9IQlfhlKzZnJuSGBWfaw3XRRdY41dK1fZn0o/3gAM1lNlzksY+xI0PfPmvWaUY9YCh
WRdin0QsDYWvHERo1ezPyeRawYSR0b32VX6mzcjM1+d+wDrZVq1LchLP1xXZjWoK+JzcN7KRnREP
8JdUDIh1/L4zB4xWuMGoal/8DSHHdAjk4FnHhvvTgKb3YVeHoHj3lGbw1NF5xMiultNselCSZ7jl
zkj6Oa7MBBFQf3/HJhEHAA+cEk4qAhBAy8m8jEyQdS8eS3mYLAM1YO3xlU4uutofw6DFLxxExUQx
eLfj71GEQUxPVWwyI6AHNyudPc3NUK9kzKcZ9VBSLJl/UMvmAGZwuN5adT6wjFgxqK+Z632GqoD4
Qy2oE9dOuMMC3ckr9e3jev2Jw0d6OoD25s6F+3FbxPPsuRCNxWBm8WucISxgAvvo0gOqQjnEh57/
VxlRV4vDjTtlj+NyZD73QJJ6+uC8w5EjgrMD15jY4LL6fv1/8RWNv11NBGPMrstjliY7MmYMy4cB
pxdHZNteDDEFriziwd+5UgdFxCzvBenqb9VlTMG3em2yw6K4XZnXFwsEJecuVWBuxOVdFMGAhI9O
tJpatgs1vMLwtxclFe9qrQepNoZmgyAnSSHliEuPUPvVQazMy39/rT3uZp7iJQlIEFTFUvhrtAUC
jEwWO/sddzXoZRHz8wbjTS/SxMxFHuLm6lffXQkyj0iIuasxZijfIe0CbnSUBbZMnlO5GMT9aWX3
NNmvd9es06sYZm/qxN0MQ8VjT7Xip6kv7TnWYSWnqSI67YbdGVRZJljUmabHzIPlD9mO3Qycy0Ml
0p9aOjctImh2FXY+vj5W2go1FIJjr6BEzsOSgs2HycTumrXU+ge7ZgDW71kHJxqcOReXG5nZzFuu
u47loFasuYKg0y/6CY2uQJDoUeBuzuZB4stLfH9FFPWCXsha+6Ni1SvGmCwt5D07cluLakeCrvUa
rexKfovCwoK3mTD6s2HbOETuSkJyWxIeMHKgEA33zKNMimxLOMbFexHM0E//OSA7SPtXTze1bjDE
HK3WxncNGlzf13umJWCDM3bR5VlwOCG/4RzzPKaTUMmVjXpzSr4mDFYQKJSeLswlEV7WbfGGfhvF
silSuKJWpmuRJujGsKBxXcLjq/uPpV1OtGKmuQo/kEGnMQ4ZXnHVme4tc8UGSjoxXf9zjxk9pE9R
kthJlnn8InF2E8QvQNB0Q/rrr/OSjryEl1VlF6Qonw9pXgEiPEa/pAeo+vKIMOnp+VUyd2PRW3vo
wH1Mx/Hsx2b3xqKo6FC9gQ02tWK7DMlZvBwVIAJvrNg0GwKgqOU/7JqpAUgD09d9t4dmkPQnOgD1
cZozeBy/jQgsxyoVussPKTPDcknWOvKTlpHHd3FawCoZEaj91+9oas+B8b6pNo/6Y51mBR83IGT8
57zss+WRWyHGpPHdyhbS31sio1NvbKtkNpBTZIx4iRowbYZmK7TxKT8V2gN9TR3JREkuoGjsQTJx
sAGrspbcgwLpJTHLHsvlyDtUOM8M+9hRziSJJwCL8aAI++aCLZt3zLo/+U1Xz4MZ0gyaIYsfEqPF
gf4TKVepaghIkssmgRq9t0yulThi6xRjZj6bs3Ljm83xZv6bM48eaUwpC1DF7H1vKg4V4K8C9Mk5
lxlDOG7DGrclEEiU0agGALqz5EUZWcA710sWu79qvF72HkUi27C/Se1vzaJgXot1Mj9jHtGsH2Fl
aedBFuyP3vG2Fn9aBmIfLMrVehFSIkFGo21k0KVZ7dBDSWbSX7waJxUuscpwEPUr44yzTuSsL+ZN
PvWclcSqiMfUYO/OuSu+LclSVwL5hDuBFcL6vmiQWiVJSJt+5OQq8rhmBH6szifR0y5XZj3Guujq
KqDqVjBGo9R5cbnCLRroDyCZyFsmJefudXp/xcStdkiAz88R64soZtm4IrQ8fuIcKu57yFybhjZ/
5bvPJ+hzL7pK82OsSdM9joqAAWk8UvTuZ/1RN4382thPHCqI5IYBSW0Z1uPzAWsXw64sIdd8cRgv
Cn7IQUzL5cpTDdC0JfNB4sa2jEDtrXsFg2Pd/IdjLdj7xyZcXg+pDamGkWIWA4A8mpHifIklbh55
31Kccs+WIQ23iDjpW/2XZ7in6AotX9M+vo+eL4vnFrZQJP0fTu/4rqjIrocLWk1XgAHFBL4aFUP9
kbEOdhvQuWHxUJsfEIoF4nvXSlF9543RCSlqF3gQUEmxiIfYQcfC5C29Xottq3L/whbnvv+A/Jc7
jN/ctcqGBLP3ny73tpbP1t4AW6LqjKs5I+/3jsX9XZDwgWWIO3lM6IWVSQ9yewTWaa4qXPu7NK9S
5v3vQyz/ZEQH172DTa2/zYPDi/kGUB8GRAdW71pCt/KhF1bVrXE4BpvmIKX1JBRaQaI9TRVfOGr5
CrnQQRu2dIqGybCinc7KJjguJvIHafWrTyYdxXhQpyNEJnqWhhVJwvNr1/0h/UECyVyvzfZry93i
Ca7/d4HBQiKdFoTw73fU32CJp3BsQ793gTvDXH5M5BPRxQQ/U10kTYB2scEG9im8qvL7sf3TTKhq
JqqWXDEqNzJFYLU9qumrDzVztGJ7P+2MwmGjkWoeZ46mu/I90maYl3DfZo9ngoIVXdbmOnD4xU9U
8I6uPS53t88q1MJACkKuySqxeuhE0iWaZP1LCj8OE/po0KPYCSFbf1H1EdufqzOJCaerxDeg9urp
6M7MORImmPDP80wXtLZmNlO6QSnxMeB5E5h1jIWEKkYgN6oSZiRu1S2vxvubiiI3grEk9KOukecN
Yp69ZZzv49jMI1MG9uQ+FJWHuc8rNBeJfVtLRoAD+7SWk0zD0JBC8wNw7xZSoaFoMjbA1ke5zEY7
pC2LUv392zhixUh2vuvW2s7NrL4TigHulbaiavpSPMNiZbl8swrgS3kx2HESLtLVmsjNmeaqjujU
hhQpgeYHPB2QEzK6c9WV23mvDGbbpJ18sv//+wpjCLrQq4NI7xsatS4v2dSJLXbociCDKnfj/aJF
h/flE+XZpbuNlqH1tl9pr/RuZm84lse0kBBM9IcSzoeWI6KjcqJg4u+Aall8BOkMSux5l/z+1Wfj
BwdRngZmS938lXcGg2l6xZ7e2uQn906/vyuG/KgbMsVocl/zBpjXk0DZBVYxzJz2PAAxQgh9tFDC
Ea+fXuuL9z71WWAeNRql6RHd5zRbG067HY+T3z+Lv+usFAeKlHYHwci0ObfLnKCBf7klT53IObnF
f/PIvQirPUFJgoFL+0Yp9oJxVqETPVRAc9oyVkRYql3WJ+3RnjNjp5Bepf7njk+VmncLSodpOwao
WX8Bhoae0kQiUpBa8hG1r7n0tzUTgXLPR8x+XGYZSoLuGA78mGi+enoNc4Ze4UitwGRpJUEBMDkH
4gCny/RJ2wwegf9AGYJ1V1IDzMu06KcFk+8m6pQqeDR4y+//qZO0OvQm85GCVVDMIe0w8ldAu3Vr
kjaC4u1AqfC19LhDc06UiIXDkHrv6759bvJmCrh+1qHkmTMLfJ00+UXChlw3sK4PVFOtN/Vg1Tvi
kaz7csJNF0AeblyYYOBRPW3kE8i0JY6t3u8tr0RRtY/Dnnf0ZGh+mxeV0GV4FSsak9kqqlCkmQ5T
JiEAViqstcoj2X3ts0oUcGTCFbnvpTeWGGsf+RSCwUskNnw7GVvq6rgFxH9z4uuubyevvhmQgtnW
Ytwl69/+6VUrpHGZkd0UkS7DBnWNFts1IEnumOdnkBT4sdFOT6HB5NMBfEznr9f6xBl3gags8hud
7bWoZ9bIdX2VbuRkToXY7nAJzzCtrJ+7OjuSNwCcm05AI92ODjTDP1efKe3NqbSN6EeFpT2lybs5
O0haABlsWzqICX3pu9R4KzdS3bdUhvgRNfJfT+6P/8WIG22U3usgvACglT/RI6npahQfP+QPTig2
vWKXg0LUw6g7PEerUKdwzGIpA3n+RS+E8T32bHvHp67qise/+Ig+3nHtsspVzB7tvSWlQ2kzF57F
UEow7/EWNC+HKJf72nos5/k620jPV6qXOF8US2QeKbh4/LB+upNM/ou8IctOUASNJPxwktoDGPnR
KNbMfgNjlU2etpwrrFsFOWEWX6MfrGFzlm2jEMriiW/sLhMhEL4gG0IQM2RXQhrLuAv2hmjicuiJ
923xdXITQkPMex4n4u7WruFGW2P1kTLx/8oBTltOmR6MxGuaCeDeZmNzv2vWO1TGTWfHXpHyKoGd
rfVV56gkKkpzoamKJmc0mD2MuvCno9bK/RAzBPkSRWTzg28AOMxwoTQtC3grr8jGloSlZlqC03yx
2/HtjHzdRDzq1nT2hf67imzxMv0uKBl5rlrKlNyh9Z3NkTgnDbAXmdT2eGom7Nbe3ivMIF4WrURe
Ud37DdjppA0jc7lHeSiBShzEki3E0qagJgIrVx32uOZwvgqnLTeMtdrswNZrHdyeHZz/uunYnaDR
2zftZajETCIObaW1TSlcMBEkr/M0+cDpB11M5UBGq3Kp1Of3Ay6lCzAXPbKMiK91yuLWJMm738CE
j2MEFSP6dLIXbdmslu52h5E8Vb1Rmc9X2WX+nEWtQEqmF7F1YrpJDq4NhWSJIoGQlaKTDZL2NCFq
+4l2URD9mTOYNqEhIf8V0hNuI1y/R+yb6X8pFkcbQtPkfSYtiI1fkXKIn0L+Aszh2Uf7P6/pl3cd
onO9aofaBIkcbRymRnVxqPoOm4DY/70hzz3JRtx6aYdO9mB6RWdJiWz5tQbb2XGyFxI7iWvGLdRC
54jfmcjld66PFGJINKjaRGugJ4n6x99/Mj9+YFNkLEpo9fE5Z00dUXHI64CvdUzzCw3yxuKiix/T
8pMFZn7TyIlIApERY+M8XQGbBEX8b5Iqd3mU+j32fI40XaBNcDnDkjnfOzLb86J6l9ek80pK0UQt
mlERdM68BeiyYUqP3XK1WSawLcGHAfFRIOJAIi82bFBYsJfrYEhXQ6Vc7PPDsK8dfxJ2Q9LlROte
zolXiL8U0ckjsByr+AWb4yL5GhtK1ZxIaAVLxqaTXOLbJXUr6oqArWqNpJtD6G6GVvnQ4/DDeB1W
w1IbjeFJ7ynmrNAbCoODn7+fMy8W/py9Q1ZP3Vs7ToPVeWQwPsoTJfG6nLigtoullAqUDaZlbptA
z+V1AtMj8SqcXqsOiDhdNJkK0azA4nAjbtKa04REjKxtW3VK/L26kuh6485drHSIfyWMDfgUC8rx
uYK8fqfRl//8Qk8wo9poNyUYNXkOt2w37IwV+RgZkm6fP0brB5FY0Xx9us47vC95mPVuCe+kxLqy
v6q3ZZahg9efEi600AJCNev7ABGaRvcGmf6Avpvhet4k01TKk/CX+KX/kQoPCBzYgTCyYl04GK3q
Ea3r+b40/XKYwDipR3i6SpTLNJV5soZCkrf8+8/0INXmioLEbpSgwBh0pm6rLxe0iYDIT6ats8bo
ET8dGrLd7tb1gQ1Mx4l1aYRz7cHSBCGg6U6UVd6nZpj6BecA68eqTZ3FzU6pMJM0Je8MgFptCtdP
6cPeyIlgxFfBMxCyIFnf/+HO3+ei/kI5GRQo5k+o9WkLfgiwzx6Lb6zM4EXITFKPJydmLM0rLvAT
dWly/mT6vJy0OX7EO1IB2XAladAzFf/hUU7fj/1bjcU0TbvGt1YoRk+YXU8Yvzh9LSlzKuMJI8z5
190zJaJb7HZsCY3vz+Em588zqHIegjOsgcL7rkZa5hm4mJ4fLbCEgHbVVeQgwhQuj81joT3JjXkA
OvzFszCKV1wdaSk60Ua1N1ILyHq+Zsh0sKEfr3JqzBLu3heWHSkoWDHL3oKaC9wxf5xem7vsH19g
oma9OpIg75P8uFm0p5CcaB9pKeZAJe1iIB7vOcG8hzOpnwc83Kz390WRL6qjV5JdWm8lBpFBYery
c9Sm+Vooz8mj7NtH4ZOrX1saotT1AAo3Rw4xvjyKpxA3LgxuqjF8sTEmxGPVgz3ZQfUuAQ5v2fFe
KRpTQhQheUKf6Pxk+lPi7W7x5ZeKR76smdRJFXbrCg9C7XW80puDnNH8u2OvBnYAxmp+GdNZV2w0
gn8mYeOj+ZFH2mWM+93VgJvR5KzspOJpRS1wD0yayGGA8VeW2QMvCqQGGxEl7r5i3DFgsxUDd7ae
s0EL6UeMI0kk5Zd+yQXosG0yuf1kRA9pIvPGDyOUI/NhvjELeDXi5Jye54tidNXH0k74+lM6n7Xe
4BhSDOAx5FKuVth/1u17b35fvyasDMeVzU90CmlAauQ8ylVfqa9n+zNJVYwlPrYpWVo+ls8w9gqH
+H98WbmKXsIMr39oh9p5uGiREaRNW4nPuUnkAPk7Nd3ySW3reC+kdaOw8y/zeCuBwKpT94I/p+9T
76icOAQaOtWI2NmP8hvdzOxiuqXlB/qxXxRtI9iahNxQqaPx93LtFNeuC8BtOXEjBhzCMfs5f2WL
FFBt86fRl8steRHlzQM9/92xcnYuvFZzpfq5svENkvdDbLzTK5jbnt79+1WoKmePai7dbGzFZKdM
2iDZdpd4G2XB49utrjLXFzQASu7XLyT1Ty3eOYjuXjW7TDXoAzYf0q5E3oRbIolr+vmvfweY/aW1
j6Q06RoIWLrqNKNK88SA5n3iaF/kwAUVBEdXLAZoiPQuNZwzOlH5q6Wja5px4/kWEFKnSdrksv4n
hwy4+1RPxiGo7SxVsatq3wTbSDZr0w1LCBpnN7oyuZXKGpFOE1hQnHebhQxGMrfAQMpX4hRk9Upa
tnnF5F529Zl6qWNW7qu1L3bf5lFCF6+TcWJiCbI6KK/+4Dny2l2zMRZAjRJzLyHnaqzGpjVO7WhY
19yOVNrdxigF3G1OPSi6oitDn8hCV+gNo1P3uZF0Uk6mROvBZxjwOspA3+bJ3CJYTfSgsFQV2UhX
bFF0BPvkYlUVyBeZa8xFJx5Q86llhLPHj3YnDHnU4mERZ7lpDYaS3At1lAmprFmDNzgusjyNvton
wWFP2takWl+JrFNNTORYCj1MEhe1HDtNi/QdNYFf+7aUwm6hB+a6ic01Bxk5fDK5FnvcmLCv7JEr
i1ML1VCSOjTc7ElQKXYSRjhnV9pPIGgUVQwpUu+OnJJTGvR/lqpHJt42eGtF0+lcjFStAR/zJaAD
dHJLRrCcxCxR4Ln0yPiggmctu2ESfWsNUNSgeqBURxc0aH0PDpHJaosbQBoU/LVK3bzNSjtmaa74
o6BrFZg5z2qvoQHH7XIk8vT45ItxskbhM/SRikqyr5v1y+MoogGjohIALfV9aYBGZk0+WeqXyeCt
+hPAK05BVgmQmOEeVblri7o3j6zjW8HzOHIR8fEB/jKWQ7q9aNExQoFACScndyN21+hx8Vs3zYxA
mbqt7E/XwTGAMdj6eMQEJG/RsT8iqypj4UDuNFvpk8ZJYAFe6rJziglgIPwyuk3Hl9TF2OrX1bTP
cyRUkPdcuOGi9nCQh6gezJ8XL5VMd6wqLiqHSvL+jvS7XSXhu0oOi4LDF6tlvWugUsceLf5RoyGl
ZNN/HqGlgBFqFTRVqDNlWnyWq4eR8FsdCjBAq8tr5apXMM5Ki7uAYXZyM80mkhLzrX2OqU2IfiHL
MpKxDkUX1PzcmgGPqLadzbqBkM0WiEfsv6lYz2Dz2nE1LsWbJowaaF97ph6Wbq2Dnwgy7PihvWUY
hKgGnXMElB4zehsYbvEQ2MeRsLj83/oZUWU7osJVm9XiOFHQxma+y+H8EXgldiun3QER5V6qmNyH
gGkhcQTUrGSs1P1EHHwtxoYKRJD3/2AaD2kl5scjzG7+FKqtbSpxq4V9NG5OBV9Xi3v2BD1azxbn
x/GdlJm1/0vfy+A1cSD+eCmMAdBR5T/OZyf40A2jUQelmkQTvK6MAQnCbO2XrCYg7zS0fFJWYDkn
R/aOTFxcOtsLPwaVccQVSSXATHu28It1ztK6A93zFobjBkYYCXSMCqyGYdzDlFGopNJeryudX/EB
HWaVb7yzi9Wd0H7himkpl1+uuGhnhGTn8HsaTdRPjUW46Frjkl3QmvwFuFeHD2gLv1Xl4EWewLci
IrOYvfnjUkXa5hOJzmLg8FDcReAAhC6pdST3OFZq5BlOSQy9LfFp8rLSVjgC0CNVvauGbfZONKOh
iDGyQwvWRDt2k8OqNQCLdockSCRXShjOoUqnhiCR4NQdyhzXpQ8CLn58LdFFbgsrRNcF4Fpvd+Do
a3Dp9fuKJKX+MnwtiVzZFo5CmCDkwSM/GaYBOrFiQhzx9+bHFpkv8COrMSwpNsQaubUMQvUbrb0M
/fe5RpJoyd50OvSrAopp3qpeoyzO/qHMA7LLj7d0d0CMAGL39b3Go1KAF7ihisDCCgJ2Sl/OoVt9
eIKeDRzgDxZZxf0jWHvyZfi2pb2Wtj4lsdWTrYVsCagMPNCoGEJZlXyIn6ZHmyobyqQNx16+Pzcs
DrSe5w0SNd1Xxxwla2Rlg+KcSZq9tIIkPe0j4La6UWsTiomQIAJ/6xhBijtxVbo2alnTou1I/7G+
x1Y4bYWVJxqMTxLcXDUSTbyn6OGcd6h1cB73ToqFn4Qv0imuxrM5uvl0U/Luu8Ah50YpmWgjjnP0
aOIjgCwiSSJnyokHmZkA3Io2sij8i1jof8Va5flFdH4ig7jB8hvtgOhU9SdS1kVUCASiCxTFoWAt
8Mbxkj027ACMnJ+a0kgogu4EJpTU4/oH5iU0w9/UqKYCHXGHDbGftJQ0hRB5/hhYeR1+B4aNnRxP
fI1jNm5BluVfPjPOy+vha6qVDlgLgxEGcgWMYy4xdZtpDauFLEU+kix26I5vQXplTEAVgMS9x30L
GFnw16Z0qQBtucKgaw0Toqnl2sXmH57BKDo877Cd9yjTup0xy0HXfQyyfa+8M9iVFYeK+6f54Y+q
DG3pgm4uMvjO+/6W47/wDzSlHEZAs2RJDfaT4zOtRd3y7LnaRNAAMvr3EE/BDd171dO2KHliZFhK
ytAJCXEvnSkPoMdarkniEHkukHxJXMl9c9IhKLWZJB/0CLGcQ1FTkW9DH8bm/oUf1TnSkvmjhdft
6tOvv14kd6PcKJu7XNByVZjSpLYQ8hEQcAduTDyVXll58sthS9ziv2PIfh2w6TNIbcqXUGQOAhKK
h+XhcPKKhQbxhjhNFSutH5XgVIM9lmrWV46bnJxamPNiyKKiWYCGwn30W4g8vrpcSLunpa4v4acz
Mjw+DoBBifhb+xCctUkuFUvrlQs36M2UHHtsoBtDeq/mcxRPymPfxKLI42x6gNhh4DOtdBSBRw/R
mL0O7bj/CQPGyff28VmriG3DxTdylErgViapdjL5GhaL/HkgcXVtz1fqfGxnSFLYflfHWf5ymBt1
jtZywOSlo5PPaqgKR+hcRCpqFJudryf9nr6XtCl5oH+rRHrr6KvfZt4Pf98MS2cqVLvTcP78KzMn
7vxR2jdYXcSala3pd3q8Aw1ygVGf6hWzmIqv/ppHtsgDoQuo4jDQNB2byWdZgVwUt0XtBgnSgtDS
nUnLRDc9wsINxAO1/IC2kt3EOyVxcQamBdNt2ixpWPZVV4lEkhtEUcS4CWuE2YxUQP33Cmq39Xbu
vW6+xxEiyq9SmDW9INhF/VMUAKipZk5Bgo9D2403wX4lo45seykLdCK6dYkKm+u6DenQX0DfQjYa
cJfK3ygeAnUCKHg3zD7L/Xxy0YFKgY5zdq35O2H1KfwYfRJTzCC0Z2jK5VSGZgFSKPsR9//kKa3Y
NX6udkwHNECr8a0S2dXryuIgSoPKub/Icu99C9YPdI4DiGEbllUJ7SH8j0C37UP0k2gR0xdIf3hO
nYJ5hsPy3I1gNlVfbiNBE73HTKfMxgMSYiJawZpK7SYYjO1qAzfRYonAP6f5UNKwgZu5+lmC8SVJ
Yqe3aCaLZTuv4yDJvqiwdbh9YggHUJ9W9hc8At7MzVnQh4B5sbW0PqDhU+IxHA8kQPib1hDtexYv
gfjB1bnWtKIe/uTJzp06P4nwVtOcy9N1W3OUdK4TiptP+GGa6C7eK4R3y7KnjHNylwuOW/Kgj8xF
uznrzZq4rZA/LlYiIO77unE52Mruqx9Ff1KQAwCnYWUl/ZOMcSN6lBuFhyRlOTBn8QRr10I4g8oD
L4hD+yrQyFlUz1IPCoc9vLV1SsngkOaeI03wM8uqbr8jY5ARHD/Q8sYJjhgPhFdwsMqUglgGfwn6
Gpg/+g30UMipLf8U7lRNcM1Do1+8vXAdb0KP4Onh9zG9Euq9l4mNG9fZt4LvQlpmIVq4hi5zfzDx
w1SGalHw9QVHH11/yFodToxW1XlyMCqItFjHB/dPX5zQNlZxdUCP9/r9mCg4AMBvteQxSKuRBTSL
b5De0GyniOYLGYjEGOAAmnIJoczssVCo9CoATwrZzP4/M1OViPBhbRJeQxmMJbZ6bKjBnxixusz2
NGnIPuL3mXYweq5KL9/bCI/Y314lOywS6l8xPdo0e1w6B+CUqe61VTeZXK5UqDggg8Jkl24okSVN
Udtwz6TTz58gUVE2tJQj1dzR+H4VBhNOS+CT/ZmLzSsFXQdOFHwahdZLZT4f9gVb/NAIvjLIABAy
IjNQBIIg1RNXo4hG0mJmzM3ebNjoAbZUuyeiFajRTfRKCDb7ujv8Qcw0LbadsRUxR/lV4brQK3TS
/2qjPr0gN5Wjk7FkbEd+4Ny03mWxKPC4Jr/mFWajYEZC8K6mv4xLzeNE19nMZAE8FmGa4Z+DGxg1
ARaHO+qR4psZSH9CApF9VJg33G3/SEThJYFOD26g/nJEVhd1/+pL5M/g0f3Drp9lccSvoroUvX4I
oujqDlC7nmxfslZDnhin0FcR8f2MdYYzErUNkdd+ExbKNzI73sc32Dmcm3/6GiPgm4OH5Py2i98S
pKTAP0l4vEBkeoq4zo52bMlONtjKw+H9Ri56sjgMX4e0vU4fgSgTHMTOaTLV00u71wdzFLXq/O71
3OMb2TjwuF1BwsZPJul7Fep/ijZIcOi4pRI2AgbV/JrBoUWIrAXCays8nF+azwZMZHwPld2T2gm4
fpNds/JV04RGe0pDHlMNk8lgP8fv7p7gHT+1hDEFp+tpK9deFBttQanPRoH/Rk0rhzPvRvakblIV
hodh+sHOFphboBBjnl6Q+WMnD2UkLW079KWz+/cG3zAypVZllJUyszG6k7vfuCCA+S5q6aYvWw+V
/GhpTTGgc3CjW90nJEgactXpQ0cSR+HCywueHagi7Q++Peoy+A0/UUMsvxbK3fqxuTkft+WA9v4t
/VhPbaeMQNCshGHx01vANEKnbOIIB5UruTEaHjggIhWZmkk3qRldRCvq7g8AOdU07GmOZpRn8ib1
025Lh0e4fq2uwbIpxUgTJwjjB9mdA/hGKlwsg5tt9Ix07CiSJBGhUPv2vLZspAc+8L8J1l9SEmhv
rzIiP3JyERR9DSy7IdnZCcR2KaXPkewNtyX5GoSrw1vlVObpHivRTTWywrGwFNPk22q6/VfYOz/o
RxoQnrqBQeRfruEqabbuo557cSq5TDDMfcobXXcOjXIFpvZ9vcspBzFAJNwmMA7wMwPaiz5egHjw
iisHRxEPbGTVB9P9uycBIQ/30WGS8NuE1+CELuRt88wEPph1hlMNrrbB9a2WlHt8WB5nPo2ZwRWG
eCtDg7Kkyl/pTNoDM+pq5T19+j0uXWFoWZR4XjI2/aIIkA25/qZWR9pwKxGqLmJV3l/WafyzNWR2
LCS2ZRoOa25HmsIvYoGZNricEHrQ1r1tL3Xhn0ppdfOxO81U4gzyDCaoAc9DeR+Svd64ayry6+oo
CY6XqjciKV350WWD1Yh90Ar64D4Gy0KO7N0TbPy38FoMycKfFa4uM2UyZgQnyxpARhwg+uRh6WnI
sE/2eLviIhD1OihxkXcFC9RNhODz4UebRQO7NDKqmt/GEpfMxGJMO8InEt4RivnIet/7JkguypSR
AIqVob+uWdYy071zm7yc6hC+gtfU2EPXD1UTbaSzGZfZuEvvvYzmPykndH22AVDWLPrhC10G24X9
bgQN2KtKbg+n6DrEHpIBtypQhmxBUMTDfQWWfhvJi4E4UQdI6NJGd+sRm4KEkdBTG3X+fmAj2O50
LTNKZBTXAUOCl0DuCpVRAMjMU153ao0jcBbOU2LkxcRICuZisRdSNeZyit6z/2jgnZPP3OamiNWa
F3Y4TniZXd+TO8/vpX36eblTy21EmRZcLVw808TMHfG05UGY+fc6QDNuY86xZupsyk8iyStdcoWz
sxHxX1mXlH9hw7Hi1Nw4K0kT+yyUOjn+phbBvM9QE6Hw5B1+56qUXCGca4PKSW2GKoL5xC7bvnE6
+c1Y3FbR2lPZe3x83QWsXi+1ERc8/TN1nCoCoOZYd/Jbm7hAv9Q0l6J5hWRz70+aYHgpuaN2qJ9v
hnV3CsA5c/LQzvCuq9aah5M/wJie4pVbXK4ctmO1QWSaXiG2HxLybVWBM209W0f+CfWUPcaAEUE+
v9JhftvvwHipSk3mm+PrYLP9HO7MUuzkr3TYZEDqcfBABCMwPQDrEoBMf4P6T8Ba2FknlvMLAq+L
Evn1qxMFJgqGU+P0Bqph0eW27h+6gEnQKmIbyaWMPn6K8Vp5EVwtnrUCZ+K+fAsLvdrxhMwKI0Qr
ISSDnV84xjvXwkkw2mHqCLBSJ+8ThTBB2QZURaCaV+nBm+Dr6xjQq8dKHSDHthniCV5cTE8EQE5Z
sryusVW8ZVI8p4cXp4uXix0CRPxDM9UbG/l9kRXaiGaCxL+jNXalqYGHaqwxwb3YxkY/A4dtVynq
W1wYc5JftfFtNHMz6F1XogRtTBA5/JWbYnQ9EtAMAB7gyWpCHI/9vsnzWMfh7vKs0SSleKd37YQi
SM/RqhmR7nep1IrjU8pCyeugsmH4SIg6G7CCQqsi+lSgX3y5CtZgXMQAZ3T7UFG04n8hYr3lBI0j
IY4e0gIJVr9v1rA3S/T3HLRAMzR3VrRKocMEXabMj/9FtW2NTi/RTSEnKjNtrxKgqaIVhfqrzR16
pYfge2p0xvtcPz9/vsR+cNpTqzBI09pAZE0r6ojkV31VhQy2WIBo+ZPyuvJRLgotcg8V+GHciQkp
JeoyuKT7fT26oeoGnRbWL2rMhgIomDk9DPimDL/Ff+xF05hWStKecRam/e7r7/IZhvudsrDDfCHo
Td1jHEv7vzkQwH1rk5rVvgHHyKpyKVTd0LvDEyYSoZ4PXH/Exgql3gc8jh0CaeFaBiSH/3h3W2KJ
cAlN02pZPuJ2e2tO2j9+tUbteOnR2pYBYDZDxYv6UbrS6ZOFqDEWOG7pppvsCQgD7Lr5pC1VYDC/
za0QoJhzCY8pS/sXJIThLa9KMbCYCwp58CUaxgxhTfkG953rtwwx6W7KUkwme2ldwJaNnFw8wsKL
xxZyf0B19PMxAWIiP92SRLju/eVxbU6CXPYG1jO9Nf2UCwaFUSmS2KsGeWhyyOENEdPPTKpTxVyU
waAMI8n/MiEdqCMxXWfuMQOcN0UjrYn8tTCOeu3V2Ase30gieO1PqkuzKhxNK3rW+yjg7M50ahkj
QTFeepOxmrVdwQDjP9VAR/lfu+Sz5XaSzl5q0SfFdgd9tHwGuxPZ7oub/dbV7xIOBS213R4zZAZZ
mbn0YaXBmBv8lQSLyuXvQXUAFWMrIhL1qBZDb2BYIs1adeIFUF8oczJ8y4+0rcRpo/oikl8CLr3x
7+PqUoLwV11asjIV0g5YR2bNUrr36IG8/91JUa6xdUtKTcb5bGh3nnpyiV/fAIt0vFvCgH32SsJs
1Bh2IPDzeatqw1ftsdPrE0uduObU0o2SOFFNZBT3JuIO46eRCPQWnn1qzdt4d+/+6sZdaEweZIpg
mCA3aIjBwi2QjzVa71jcFPcJReQdTHkF9NhIsONOUFFTvPS+XysEGPwihiAgOXBy1HMJJSzBH9bb
cfl9tPcme2M0GF0FlRad8uY/Iz41A3fh0Zii62/nd9rrXt4LFLHEs4SWyv/JdsbYqK99+YATxbjE
5zfM9dW0HLx5hXM99M6S72BWGBfrQ+i0RdxRKFwrRcQht0exVgm3Qv4G7i82kM0lBFmK0Uh91Uf+
0uKDnQPPd35NBzNe6xF+jvGsj2QwbF0d6R5VpXFMzelkBGMZqMpUL+vBioOPJyjWiihfQoq0m71s
I6j1PDzqgG5ONYivhBfIz4WGvL4fJxj6MVNYRmfMij22eEB9ttJ1zHFQNnEReTuhOZxJbW8FuphC
ptRG6bn/mxy+6XwRwWPJxuMHpJM/m5T7o7zEYkFjntylfmHK6357aV8P7t82wahqSxxcWGIgCuiN
G6HEBfg1zIrK4lr67ScMe8nEvxKQ3Gik6sSha55ZI3iApxdP3C6S2s2Oj7fMW7gOVp96Lh6YkwvY
q7dKUWd3XX5uHmx4/c13KAaTnFeRDV0mAPx0gt4fzxNF3oRoukpPIwHW3cwVNPzrjBB5xImu9XoX
MbLje6G0Tp/ercSKffd3oz1ju8GS8JquxPo6p1S2rwEJq29h+jDAfKjL2ZSlWKgLWhlY58m/1qVl
cffzayM6hBu9N7W+XbttXjg2xJOCl2nyvAH3THnzqfahkCdPZOm8F7jDfNzxNf+6zjiR44ai0myt
MFuEt8rsdvQf8reQdtoaoabG7DGBmg+pakF1WL7p2+nAYtYCRDGPwYM1Bs4TUl+DGbKz7DGoXJXh
Vi8PtBFbK6K4x7Uly53A7Lo73skVjpUxd6AsgOy/b4MFdeVHSZhH4Av/LKW67usKJYsNv0rw7ECI
59hOTJAoMJGeg2XOZNCqRcNAA1EKszaFub7ZLrSoeqm0YGbAK5c314darqp/e8dp32dqr1uN/ouS
fwdhq7NgeCQYhIgO2Uh7+KUWvVOMJOeBd92UbaR2uInV6ZdvcnwevZILwfMuYPrk+QPIGaE/n7Ul
406LX02eVw0WbyYZf/pVQFdVmMioaazxd2SlsEAPtakOZdDyHMKCua0f5+kdNz4sS2mJgx3dk/L9
ohqb9Hj87U9dY+yueVVe1dv3OFKWMuq1W+pqNvB3JqujOCL9EjJ5d5qNgymAc7Bbvtat9rFaNZiP
iqCuFYe1tkbT6qV43LgAOjppxBdjB1at7hEQuqo24JgWHDUdZK4OVU3A0KXyhbQw2yFcK8gfoFoN
hlUtsZqBOq1A6CTil7AvfSNhzvC6DPs0bpd/xAeZ0A0W0Dfg0yIUyBKJ224sLJygRW2sKV/Vm/eu
uzCjOtQGW9FQQR4yWfm9cWeMSqoLk62iwecrFKOJ2AOhIxb8JvCnwSo6qJX/jBz0hiO5D/Q5F5Qa
/BvZMBm3T6tIqYp5TOrBXWqicuV/TDRzierTBu4M6wdTnCg2dThShaslivTnRX8HynamJLR2SYlU
ONqmYJOSdpKbi4LoD7uaAwDDrarCl5VYpGcM922lOwITND+qF0XHs1ATDoGFYyxON8fi7JkBkC/9
F+3sRNzBrULP6ZVFrsKNHxsT42tR2qnB1MX+E6MDZHrfa3VtcxQnFqUtRhtSvOTxgUWe/0ufvrFB
s029awy/ecF6fcM4Izy3ZjVgV2toUMmE8HtIYuKpn1rc3BLV8gMAxbrC4KWlCnZk4dCSqLj/bCsJ
WH7OQokQPcfG2E3oGN6UwOtpmHbJJOAGOZlbBo/WpOSuhWHa2BaDuy81BI2VRvSEbroPPvPSFQi2
aCYqzI73KdsS9NcwHMw7GEchFuXv5s/iL/KL+LZxum3vLOsyKhh8F6Yf2bhtQNo7BmuuXXgmeXm7
s+qR4cfpcoN8ctZYMyKmFL98AVb4NKPcWf/YWlYp1RymtceVojGRevWm2yI/p/xMQrbwmvWtV+/u
1mQ4qbD+WnI5iBsRUBYz4mCzlh/KngN/MH74qr//S3hOKl768Oh2xeAzfrFe7kzj6F6yHRAvdE9M
TXRyVUvecT3VZcy1NAktR/xSkMhpRmhzyfB3h36BY+h2Q5V8jlbKJgYVzj9SIUkUWESX1si4PGZs
AzXaCCSsDdUuF2ztH6pqiXguTNFZpkNdwKazaclWOs1vHnQMeZmwYOgA/fgMrzpeGdkY9dF5m2yM
Jrd/nuL051ur1d5v7Bg19oh05UcXEF3l7Y3/cGbIMfPFcdQZul0DEZl0DefG1aEawMLUEHqRsbLh
QwmIs/mvAqT3dp01ZNJ9zHVvPm6OLV+m3+gdLq/5jDoocEEhOnMyOTB+mgzesaE9gH7vLPJOCXtw
dlVPt7Ju40ktkMjaV0Sj33mkzJHrKJZmFTkRSrCTP89IyEx/YejQeqaAxwRBI+nSO6z+XxvKLwbH
WMXpaIKneZns6ZQY10qsxAc7hkI4d0260blFPQEZSmVmyXcJtOYh1otPXtAsr1QWV23SUgv7V9mI
2E6KJXMu+kXOCaqdBd8ZUOGPTjiMTUzdO/JJ8DDWDPImYvAuGNXztRGuhGK+Vq8FO2IdwY+UFaaB
jBULRURLPtBiriSQHRH8WKPuSQgN2udUYaLbgo6HX+fBJ8xcT1HA0z7SS0vTszaz6IGc4P7H8Ygc
ZBEbi63A87zZgEeKUnTO50h5XVP+zcH2CwoUZ8h3rxE/AycWepSFA3TvsDf1Dgj7tJPmSNPbAo27
Zjy05rJGVLnb4uv7Xo+1DWGBjjif46uc1fLg++cwatE7J/kWF58fGVYpZQs3xJSVXqMLCkEMwN5k
EqCMk1EsL5xWunUQjGypKDf1qi4AOz3HCVaEOqF3fARgrx34MZWG3KvlgyGLjdLoScqWLNVzjcWd
GMurbr2JLDKKtdLuXK8hNiDrhtOVyijVwRrgpbseLuDr0R4vZnn5hj3ODnT7RoOZH+00WPyc2OOR
dS6yrwih9tcF/lSjkNVFQpPByRtvLlTraMv1ZcSqKJh5ShpdQ+GScXLemgKDKKAR6wkhEHibnqA7
PnRFabVg6eDb91vPGO95SOz+6wQpS+v31r+8i2d0+rMJnJZ+nxsJvtm7QJPZ7hL8Mu6mSNeAOusM
0mkHH572zxbhSp8FLoXNNJtEz/YLcLSGq8PcnhgXN2KTIX8/GaqEVj7okPBq8bRF6XwfgjD9EDX4
pDptSlqcVdBom1i6WO2RuBPVvr2c5q3P+UwI2GZzZPnt4d54N5HVuZUd0VRjX9fPvwjTqS1OuYPz
ORBMixUDNfT/lmUXaxvV5WzRnP6+bYu9FQSB+10aqMoqKNqJNguuF5kkLtnJhZHrPlJk1TAgUyqZ
nREhSss9sCt6ZEsQZoo42vw1AKxxLRr+U+5j69WLI1iZaGc3Jq8mUDNUwXWeUF6oTo9xI0WJIvS5
Ohx73LGyRI1gvPvcT2iCxO8AMAoc2tUYTjDO3okDWg76NKcuR6e5g/ffIs1YxXURoeUdyuCrE4gf
IsPa0OwyGa7YoCwnlkC9gd9+ZzhoHJw396nCAH8aM7rQVDvatX7fRIW1EAYpfdfH6tyaxH5j3TgV
tS6TF/ewgDfJ02o1I21FGtkYAreore3ZgKCRSCzGFU/N7Pp96m/IzAmY8xZIY82N5FNe5S0stP/e
ZCyolRouWNRFag/gR5rJFhgi72xT1B2xtgXKOQeMCA1ZJQeYwn8UbaEsyclUjN06UPA0Pz4Zh6PN
aW/yH1KYEIwKFsG86R2aiR3U/d/Sv+50XDIJShEY2WQNGveLUjF54h3BVTN4pQyM14lMqkw+VAnq
xYS9C2dL8sxMqgRkTM/s4+SqDxySCIMoI4WRCsmfmquFfGtxMp2K7GkFc3Yrrx2Dh5YzUxg/P+zO
YJuDWSPWR0sTPNKJlQnBruaFaE0T2xpsxb/sEhTO4rEfocIr9rg8sQ16d4jPeR9N8WhuPAM97NW/
QXYn2QnnlezlsjriW7m3q+np7Q8ui1u3KTMUDxHoqORKZMsTF7iYAzQXQduqN+b6lEr8alBM/ifj
l5X2EsR0Oq9eAbnA/oM/ORDRU3owu5Y6COUMx9ko9/fAdVGfimaznGcy8uTzS8eDO6PTIVT3c1j8
Z3vAFQlm5EyME3zZ1EbPyEAx+wQpl/77/wlDD/OWFjUAVM+4DtJ7VEXbJcyi1a8noQfphk7Y9uY4
VO+iJZqtotrmMIdE5+KWPYkpBDrHjOjg7zjgnMSwSgeA15IGKi3dgd8R53RhyBPAvFfd1RyJKJzq
hA1mPb7A/GSJf0h+ja174x+GF8jk+FUpH8A3RVgoclRCNQieQR2rFyn5apnsvO+45uPepMK2/tNW
UpRvWBgDXYxqS7kz+TUIZzL69ZZ3mDBM67ztaM7lxJfCVBllL5gfa77aYPojW9Y1CREayBJwfLE7
WrvGF4VD8kUSHeUWuaEC17D28uaJ9iWJfRdbZSSLm//PizVwpU72Y3ssmnmaMPuzV+dJJD5wK91J
yiFXnnh1iWk7vCF5NZUspI3M+GPbH0edWBJJnEOpNPcub8QQPo52ywIt3z2jyBJTSZ1vFLazPdR3
XVn/P7I0kw2HkuJNpLz3Oj5RYVFu8KFdx7R4v1DwdAgnxFWgO0qykR9bmcfslL8gZGwatp8/RUpg
MUMnCfE1pfVKPWf+msshIpCLZ/BRzzeKiZU6a0Aon6vQftPVoRGGbAG0hCjmzfo+6jFcfWqizzpc
nlBALrt4NyyKgHHuZJ1iIAj52xd8jt5pG6fcs1BsyXK52CvOuYOF4JF5fpsCwOAN76H0AALKDKhM
oYeHMbUyzDP9Ft9PSssoJhJz87epxwtbX6vYKRrqZfgXunG9i5fxQF28e6CnhBL0VertjKfU66O3
hBTnEeP4DnlOQ28tv5tQM/2ZsiTjPeSpNr74ji/hXsvpQg6L6aC4RabknwDz4j8+DW1GZ3W5rAzX
qTaseWjI26McB1utO/7ks0MlGg94tMn+tPel2EYzn01Vmu/InfJOqUGBmVE3aVp9mLSlJlblYhCD
VLlHPw/5nF82Xra//F6oZPh3MpnDGn0ywoYjlXWnkWbTFoWtsYoP3/Bd9Sj5TGYCrMEysbQZikUx
m5BNWsHPrTxI1vyBrgKqg33glBSZk0kzBMp/2HWLkCH0nyVvbTF8s7Rw/eXRXmCwB8t65TMv0+x2
UXyWbqiW0NNs3vIy2A6RwCtMFOGsUiJg3wSYfYTcMFMhUx1UGOyQ5W1tJ8NfPdhR6VTFVBnMFBq+
SLisiV0HC91amobYvYIw1Ha4HhBqfycN61sE+T+lQQnU1JI8ywPm0iUiZc8GBkLixumxllzgRIfr
0C3yzOe9JFGX+n9bhGa33THMc1Vpx2lR++1V3FZCajSR4TIRIFrHNka5tkAabzCdiizqtrw3pmov
5C0+JCEt3nU4qjdDI+ZFNOzlqo+cH5enO2HUaCbKxYuns1AEax28D0Jk2m+euc+LYHh8tVet//NO
K1SMffh5AOEg1f4NO6EIhCjwZB7fMNdiyDc9im8FcsIKhOaflEsEA7cqcStUJ1uYif0zV2WyA6c3
yfYJsgeQiMmI2XSlafSoDG1QgE4mBJRb+LlUJKvmEfbp8ERFnQEZl86kTXF/DD36FENCkeEqEmSO
1SZyOPBAWhSku4TWPrO68uPkRNN4D9niugf3dBGmLaPpWUouvYZdcuCTM4lozDB+AjYhhQgU5BBI
Hji7PRN5EXUch8EPC0Yw5JJkKpCtwSB+luH/LjGeL5K8UqnYmR1iMzf8rpuivDa3xQ8mDt1ibe7U
AV6JF/XO/0V4yg0BNpvDY266bxlBM+p+boVu1pxT6ZRpYO4XM2WH2D0c+fRZMfmkToh9YA1eMXU+
SZ8IJeUlYu0Dm+J+KI8YjECQaX+yXg0YBg1u1hLJQDK8BnRiw0KXNNI/gb2VaIpHJpvgdgvWBnJF
j1io4jGzSQRhPwSWcV5EMVIGpo1a8LsxMPZd4z7s0v7df62Dg1Ww2BpfX2/S7FLRU9rC4rBWjqwE
rtVNYUVTCp/UzY0FYL9LR5Y9H9HGjQKBpynIDGfiUsgL/QIpMolzlmg18Nmc+qn4OxB+5kV2rjJM
67HJJclZZiVbI0FRtJcbmFMAyaTznIlVuul2F8jcSqZw2Esg91y9ubvMXavKueUZaUz//tYxdJf5
C5oir7lI6NcbUb6UXOBCvZeRrBSfLRszHJd/9/7jGSNG6l7sHEWHV4b0kBGADvltP6cYptRaPL+e
37N9OMQp0nbZnSkydy6yPdM7vWMXC9oGYGUvhSMIRoPnAFZl1ZfiykKeRZpNvafpiHkatC7hBC8w
6KUUER7nBGsCxZiIcte20hbDYzc/eEFHi9A50rBMiaD7/EyRzvcQo7pgICNp4ACdDuRoQ5/obWLx
rmkB7ZRv/eca0nG45COIFlxoTyv83MK3FUfi8NcavLN+/1vDZtwtZi2I39RKe18h6LAIlovXNRS3
2h+BEbE9SGi4RM63brWwRuStWfc4gHRA3JMsicvv2aD4HUdDQWHtAHBAANvbMzEKQXDdwKUj6h/V
Cy7YyAK7I3Ph7d1hfP0AfLiHkDuCafB5BzBmilUhXsq+2cXIbvDkhJYC/ntmFnhz83LEKyebzaVk
WPqAmet0Mo5CVWxswucQ6d3dS5YuzAJ5Nwxy9HlXU4jjFSrFl7MtB0JaMjQFyn6nH3Xs+F0gepCb
S50h5BZdGME9/khTjqRjUwMQsk1MVjaGabcHwHey35EF9W0GvbKqlYBiJsDNBNDWJf796yr3iiUz
9tZCY3ghHMwcinBoVvlXv3o+2YCieUX0iPHz9rp4VcArh2aHKn8ROwL+ZWkOjS9aEdaahQtzHZ7U
HchNRfesFD4GCI4b7CEURe9f6LQ4GGoegQXATT/dlxO7FJLUvvJP80jjBUA8387dEMT5CvVVlBqi
PaQycZgoDBJuKR/X3M7HPm8Hv8YL5Nhg2eD716448yxLIu/qERYJmEXJsPzvyjC5z9Bkh6KaqO/x
ZTdhUnn3xra6WEfqEBY4H/H5MVs46uz1yJM4bHeF0hWinqs551DgBvQHXpZnNgEZdsk9uFhKcOnD
GHFfmmzsS/c8qcV3+B5PUNKX5c8r7uhEVGh9cJ1TuaAfWkKRWRQe+vIzeIWXrtKUtzadKAE4BPEH
2zQYtNWU2gg05rvIfCBVlkyVRNI0lULhMTLoP6q3dmsiEOdbaFHuBN6SnySX35KDo68i2KxTKs2I
CypIWtDM9+nLAbuFg9BozuO8nr637n1WVvaDn9l71PiH4L0MGzCsG4rVQ8reK5yfDn6ZBa4Bm/+5
8r2tOvR32ZIRcHAtA3JTwvFZXLIKXpMiyJVKDciBjpvgHbPVYX0VqiSBPh7TTfqqkH0XrCBX2HWw
zSKRuV25kp4ZPxK1jNROWabtOzJyTn23YfY2uhoowTzhsLvgy3SERnUuIqkm82hgzmI7T1WaTqS5
9VfVuvBKPMwtR/lThKjypjDCmRiT8BuwC5fkVi7+RgT+P2jogve2u5uiDKEWrP5P+3hiyYuWV0ng
YYXPpkxdNI0LN5X90u9dDGcNxrawNwDSgcUtoCHOALeWdl6eFTnK+iKzIi6TpiNGppQ75zO7UF4+
CmtUYDY/4vkInHkt3X1WT7SVynneCqYSBsJMFhLp2Vy1G9G8pwbxsyak6/SUbiOad3ngbhap+j3z
I+A8jxq3Q28s0L7SnOH0VPDqioszHNOjVcKjMF3RUtjH+BzoBeUZGB1YzhihHKF04O71ep570oDR
jLXOTPBa4d+/iLlWlcwZVGrTe5KggOUPdrcW89SzpMXFJ2mstXvIOo8ceYqEg52TcIilBJ1QDaek
B6AlcyxIn0r66Z4sI4dgeZl+Ghp3z+RF39n9AszVzlFibJ/iWBkhB4CHemApMFe9XRUw+fai6y24
SwsApFSt5AfDo10oFasd8rHDalMJ7cmOcN9btfVwrotx9fDJOWDOAECwj2s4OiQVhuqRmF1Q+UMS
sbCIPUF5iUvGMGJEAjN1QK+nwvEyde06b3ETsHnjQHqpnb7wnBSBB9ihk556bm2CLGvUJv3QifIa
MjRvWr1bvA3nFl+H9pqlQTdyPEB+mPha5lnsGi4Bgc9cFv/RaSI9m4rGrGRgMoQIxysbR3yzzjAD
m/yaVBAPznhAA8IwipshXfkX5PpddhiznK6h3yVHj8RqygZKd0Vn7tReUhIxUxk6NQdXJp4nHO4a
ZDjY2jvZW86kZjEUHJ9G9k+q3vQGwN8s/53egCDpvm2FTffNWYZPIt8xAKjD/LNhSuEDf1EptOKt
zKGEOz28GhT2QdMHSRu++kGVWJJ0FPc7Brn56Kaq14Z3n2zEo1zciwU4/pNIV9zwZX0P5cdaK4pO
Wm8fvOIZ/hyx6aEFNLH0RvPeLasjqX7gUjj/T2FtiAiofqNBQ2a10yJiVTV9110LQTD3tZ7eNFHu
fbIGel1e1qKFIWHH+3qspGccbrxquRWzXIolLpGbPB74sv15Es6iQSmYLz6ydXz4yHG9WIcBKLln
qDB7Dge+D4IX2sXzkYoDcc9xf9oMVDpQCPvNLSKChHyQQtAMAtv1sO+AFXWqYdlXV8PIn31Doo8f
NnpnvE8zZbO7cuM8dtvjaMRccpypnt30PUKSEo409TYgL5t17PpzFX2IWjFgoI5X72zrP7f3IVF7
WlUMvf8euIdp7i/QBuIFj/IPfdfUt/6RaDbh9Ebdnd5N7GwHwBfWITqG6crVqssBcPj4o+3N6s1I
bWqUg5wZI9YPZi8RKaW8EpyRJifkuA583ymZBLphncLvN6IfMH1SOjyplbLXdhXf643Ju5cf6u7c
tC7mJQqHJJkMhYME/OflsmN8qkTFiriPIEuS9pk56p0rkHvJza5VTSeG10zY4oIUIIfaZdU+CgK5
UDt6A5K3ynwV1oN7I3Mgbu9jRudr8EAxPrNzdoQ+2StmddKNboDxuPrKD+DkQYwxm8uT0JEdXHME
XhI8b3UBMQsObEujwAojOTljfc8aZLYnElFMZ4BT9TpxSYEYqWojKdgXeFL/Inu9En6nftvwI79n
Yc8siuZ/K/JzLdZjWU/pou7Pc1xA9/eg28ROrs83owm7TcZKGAO/PwcurMSwtjzRqy9eqq2g4/FE
KGwhqnciW+NDR7qIIb1OIwiD5LWODR91kjrRiW71THEGkgPqIWfi5JG+JJnoHIzsseY/qiygvyfT
iIvfTGIH01hgrhWxL9FWZjEJQg784GuqC2LPpnUfO7k35sBa6A3E/co6HDbDRq1ccGQX03ymBTPr
7LAigVueEKunpzzqjC+aQ4O5uplOoolK8ZQvGpkCCAeI4cyHKzt1IJ17zWBMbqoQFDyZrb7pz3LH
50t/Mn2BoXMc7wTXiIE/WR4WHQbQOz1GidCND5lg0ANv9POUkP9VbSVnVirpTsppIO+h7irx0c/B
vBpJ+pkFGTtHxP1CnQy5pVwj6Er02fEY0DeS8PpkeCqaILnVUri39r4sE3o5jdxJwtH3Ehg75DTz
FR6AlwzeO9Arnk6f5X38sokxmcsj2l8HZg/KDlVsPrq4FdNlKWJ8UuFfL8lXHJZs3d7QG98JDruH
d4YxOL5AV3SpmJLWN8Ic1avSiVqEQ1+TKYSgBKxhWqB4ffKVXWdeizeQ56kRNDr9T4EPEQfox17C
vp8o+VCY3UnWo+4c8fr97G65Si4KpN+fme7j0ZsIP8xq+teaGgCWqYwSNRxsH50p7DI86rqEB/Vt
5/DAiPN7J9ohRDS+nXuI2nZ+/fnMR1MG1wGYAfEnpIuA3eK73pYtwXpL5WfPL32tDsNHO6x3XwUy
h58a0wTTv0792YCHadXgeKwdQremPwrF2n6m3g0TyLmdkrNqvKYWSZLOOCcsjNFTeqWNkIk6eGT1
JHhruoay2k9JfDD2JCjhOe9e7Y1iHRy/iHBJzyyD5z0pCkauOjdk9OoDw5lhky28xq0EBMx40eEb
j65LW5GIdm06U5QmbhUGB+ZdkDbIOyh4gmykmFOXWGfJNGt+++W3vB0zvv/MY7k8VWFI81xiZDjD
ooyiH7M7rK/by/RTMqyrv9RVfJpYbjzTf2O3qbc2NNpOmntHFVioQ5X0PbKEj0vLXoZ7yTgOsZ7d
eLKiUJkUq6G6AW9kcjumEBcLW3TakKrqUQVqASyW6vSfzgnC8oWlt1MfuLramLBQfdpoS6Z7JCxj
1uGpotvSP+WN41xstqraMMWaIIIBSZ39TqRzcn631U8tp/Xde89osmBbZ5PwRC8bBx4b9SXip4Oq
3a8ryk5WmRfrUXO7K2DiAerCiLrSOF8mefv0Y1ekepgiQJ9y6545y9eK371xLeFCUFAckMgqvTLD
tTvpmADzcQyjhjTr3ICuUTseOMdDh/xbnxRFph8w0urnGtmjRlOnQuYVD4YAZoMPEZXGpeIHXz1N
gdWlZZMWzVhK6dqNSzfPB9NEvJOTCrZqvC6JRH9r7EYTERxXFrBeZJHRI+LZgoLqL7iykIga00b7
dibhPpOj0Z41xYY7Y6PSpAa1AuBaiAFqiL2gTUoQzpfpeU5Le3ot12uIqp5NJixcL+rQMOkt3xy3
H/g7BAgUYpc2ZNA+uXMZnDFgHTAqqOjYIkNLUXV9R7WGnCRM5CxblypoUDoSHbUPgh1wjePXqNfe
sVch/efa2TVNYfhES0hfxvYZ/lX2oWqL6FjSVUVSi9vxpwvBClJ2UY3sT0bbMF87vYcMuaPT4bXw
Sxk5IIdPjYnUv4alM7B2yVEBkq9BM4Vdk0ulOab99tJuUs5hg4NCERwQVaMPs3UQV84CK27HThay
JYrSmxXq3y57abUT4JmcR7NmUUJpRMd5A9q6rYTxDVkEMdtbWybwVtmKgobtmOOH9OID9DItVefL
z5oEl/hNu+TqPnkrINx/inerz990CfykriNx9DgfQ37m9+oy1lWg57Y9uSfOESMkZgu37OT+YWWD
kwK/d/Z3pNByoziqeJYrn8sS9Bsj9MvWRmvn48hAbLbvEYZjRNcdRalipJygfJ506ToiLEHz514T
LMGM+lqKCx6KhU5zNV/J6zgepqQcySQBWVcXG5Z3479mnsJ5rg62Lt4D8qg3vyFDC4VECcdtQEEI
Y21RU0ywVae13MoqgHjpvCEXOMLgoydO7MTA27MLgpVcBFa8QaxUy0gehc0dVfVpRHf8OC9daWyK
+ywCKWrPNZVKR/+i5Lvj39dTFj7XQ7ttAQ2HDkurWYtFAy4MUiNwy0tW8XIePGk0Lne4fwVcxyMN
FyV3VR0WUjis2SS6mRSehMaorzbaRlijyD4svoS0pbOZH/HZtQiVKN6qlYEJIJQn4yU8Ua4AoPag
38oF5wWJ4as5lX/cW88nDnqzC7wlEHFOvzappQXEDqc7ksrK4enth2L3bxFIG9pQ/5EFrOcCsveg
U1cGJZcFKeARuN9cl2mhsbafvxmriw50k70gjDjLtkzxlrhVve+wMpQii2VkUvsE5lLdwOtlWT9S
L4dnSaPzpMWle5jAszjw4/mEGuRorWzr6Qo7PgijuHBV3n6sNl0p3zsT9xfbT5g8fA57l9/kmIV+
8r4fSqAE8rKH+FZoni/TgIquTzVDDt8j7YF4OKKOvC2gutmEZcHBGwQsoCU5kYCTA6doD7niQ3gs
5pgKFD+wV0f90V9iEURoJRLABc+TTUNHfefuuzhuFUdg7+5fqwJQ13mUCoenqUidCqoM7KMfaVvD
VJOci90Fc+Ci5wCLdnEMdxJ7cfxUEMf52s7RsPA9Do6jiUl6MlNrZz9GpM0NUD+DTAEPW+FE/BhQ
jlddXQR2zdk80lFcgp5SIVXxEo1KAxOoLCa+QOkxh8nQBUnn0DqUvhF/9Intle/Fw8DEVXA1jsU/
REyCPTjkt93A+v92/qMeibeo3V9Pcx7C1hlmnlXA7+mhnHZ1p0L1PYAoizkmWu+DKNeNJso5UF9I
RauZrSrrD69+kKAWNs41u39lMXb1Ozj5Gkn98hNbb0AprZQkk1BlQNowiKDekrELktn3BqH1Tih9
jCxZJG4sf8xZKoTbMoDzqEjEx5DApDwWFzoZqKCIhklxBofRy0N/PV0FtjkNshZIR6CgOUkFbEIV
q3yCn6rwyxq1XdgTO/mPlKao/C+kAWnUfbaS1iXgALcXCPP7DMn2O4EfDXFobdfsNGrmvl2vGca0
pbgw/jwEqWMweGBbD2iHD3yFQwOD0gsjy9gaH/jeY5vT1qpv+huOiRdpIFdheVFmcerBMGekU3Xk
mpUA/mHDBuBRy/04awbyi3LFWJ7Ob9rjSpm0UqBT5Nnw/Yy0PYOS5t5eVXVwmgkZIgRctS6oDvLm
O5w0WWbSXdHpUGceh7qsC7RuPwgKIHivfixKrxfND/rRvVpkzfp8HIIV4FZN9g/FGdFFX0XY8uJi
yRsV5AYyovvoi4BGWonQ6h79JvY11KmRIJfge+8/6zFsw2Nj17NiPfworBfXnQoq9H0UfQzMXwHa
8Vv/fDNdfJFsdTe/YMcbpYOa34R88ktKBVixdwoG9mrDQ4ALnxVKOebFeX7q6X+WddzoaOVIr5Wx
MWZWrY3/1STGbxKUtWWSAOoEc7KxwVeFLFwnUEdll2RZzerccEaAPXc8QFERdRLZsdiDiLyd04+c
LW5AonR0FvNJADKqsy9EA1ro2ccvInfUofJAQjROI3aAyUZSYsvexbwzmOdpEu+IFK9WwrH2dHl6
Ktgdl8D0y4cfzdRJezEM9HPwAxh+SCXhcbVLZUGxXoAhALi+bbYj2U+bJk/HiMiEs/2n6MIGItPY
i2pqwI46mPYKFoJ7yhp71OdrAzOb9fU7sMsAC/icOdNm3wHTuyZ+BJ0wxQjHDZUJ7VXu2yzXnzC7
fCTNcNYsapANfSBjqkUSB2M3Jl3cV4DoTbo7HwJ6JopYAHMTTEYCyKYOet2CwIdbXi9Hivfkt07U
S/MjJjc82YgoqZYXH3YyZYHLI2mtHXUybaEJiFc+8YThoLEZNYVQSJ5nO3qoLPylvy1CTf/j2+n6
lx5geW9KhovI3Xhh0ZSHiI5ZvbeA+owmOcSF11uy3sOAQp2OioE4tHYLWR9eHlaXHMdXEClb8+Lo
do/fKn3y2ykbJoddiaNSVFR2VUu8102ajya/r3HIb8wSGJbn5jI8DG35sU6I0Vk4pOIxXn6zCANF
eCfRt7UmXFiBsjUDqmbNvUDupfDptKWMWiZ82eLENr97uiBq4sb39yGpk5xzWbMFXkFyQwytlAN0
hFQ1IMip6cMd4q3UjWSCJWiD/YGD1rJk7bj0IxR7DpBhQgFHtHIZZ87g78SIK2BHI/VtXLAg5qZ8
m787HJ3EdAQz3aUxUzNAqajkojqi8PdNoqxaawSX/60OdwjiWfE/F85Rkz0MPWEK+Cvnhdi+ZbAS
gpnZIJw0VtzUVLyJtoLn9YoM++9fHeKEyHtrivDNWHnKbqc+ItX9/ay5zxIYtBG36kwyKVlFRs3P
N+6cEztF+efJKJsfKIBpkWXIiPb/7Z2viFMZNdoqGQ11GcKttVAxobueD7kGrlytzzLQGExUkFsO
qi34M6HrzW32k0jndY3w7HZmBNaGEH5Oct1ldqH2OYkHkGysJUp4jlT95+jsRI2flecC5pLMzFks
Zc6r1OyBkfBdaATUAOxUnl+zEw05nThDHjVx7/zfEPI4qh1o+ZvkxoSep6yexKBSeGGoHh4jc/AI
tcfxS4FnF+KgwjqEWB4byzc/2+t7DDXhHKe2Gz3uOT9Hp6BXZvZFuLsFzaCt1h63ud1EXb/PUl9d
0bdklQAD7kNJwrSqIleP26NXfpDTncW3oEwbh0jfmrnW78k7mvkTyTrNqK+/Nc5P0ey70x8ASNg4
Cc2EHuFFWBJQFwF6jmIQ0kYQure166+KfFPWqRX+4/cB4M9uhsu5kx8vvZlWljQ/EnHjBT1vkzJq
sSP1oUX8dnvGrROGSXFoNQohriSOyD9Dr3tKaAeABjpOZQBOr/LgsLDnKPDhDRtJos4NbHCBMgKy
TJ/x28AVXYv1Ya/lLwylmRuWs0l/ZJ85UVdnCz8GYfM8DvXdqeXTGwvHq5ZNMeHlfRLwXiyGFSqu
Crb3zCoM8ASAHCcxq2vNowlSTiD0CABy5jJXyDmNWXHoqKv1o5zcAzMVlz2MVyWYhuPAFSQL/q3u
hsRSNH+/HWgY2dKBphx+xFutLnpWwfg2noBnP2dNQeMtjF4JzLE/U0IhR1kowTi3zMzlnNWKoadX
KRGmPV21QMkTNpCCkZeevKJ/+dDicnurExn2OYlmpDZ5touasU3ByeF/1xNzdmEXn33V0sZSiDt1
vG/uWCg4G0kuxdzNTGuXainsXuhFnMw0YxPkXcWW9zUoboxisxbNsvF+yUR0FbB3Kap0//rXtqM6
oSW99lgJNTg/1mnqhTuFa1e/YRLD/FMgjxAvmmJwqZaFIM8Fs3GHNE8vpD8nqLkIrVOa2NdW7rEM
rm1w/LnmeIkeoZHppVQ09gD4rpdBZMM0TT+0fN+paX9dfJhEr8gPCyrvy9fFQcK4q5t8bZ0YbO1O
o01Adh6d9L4AxUjWzYy4kt5+XnuYHmgRvWukoEys8sF78JfzWI6S39Mm7d2t6PjDCePMKBNrdwEP
77VXn2P9hBvsTL9SVksA0ciTtbSpYmNwfsesKyaeijn+yBsiwXqyKkq1U3/phczBZ3jiQUf6Y/bP
5qW+Ap+cKfinGsQqjrWQ6pIk19A8BeNWTdmucBPp0y37Efzdkjuwipz/jBtjG19LDTHtwjemgYWE
4NDx8LfY2Y78LRm6PsQtdurkl+MN96xqRRZkNiREX9Sy37KVez0QLAbAt+vbhihY8U8ICjUGB17d
Gp5IDQZWWZs4CLKT1RgOVdWznsHGOM7LPHu1U4twE2ecJi57bmTBNemu2UHEpoOHDkVprKyzVnzy
HJKYvc6m9ZEaku3XvLYIAqwUD8gcDelzkXTA6Jsk4VjGK9yfGW2IoqFIdVZFm95SHnXhkVAjfNcU
9/ByJkdDctEZ+wvH/j0n3WACRUWCU7uUf+lBmxiE9s3wZIHKqK0Y60NGkAxhfBo4ceHV6wv5Ctsx
ULSo/cfvqk8vhY3iD0o6qqeN3ewD5g3W8lFvlHjye/6sE44jCG4M/o0kZ3h/u98soa54xAGupYPi
QeZ44PvfYVJEajoSNKCFL9QdNHiPqeQKltm2j/0ts3db9SRVFjsxeLVjGya7tg4vZeTDpGeoeRdn
MxVx1cfjBTe5NxM7bV09XP7kF9vt8pUGAxL9uoT39OCFWy02gt71v4bG8720j4bxfOadUjwSqq+h
kW2N4TNXmTCRM23VFGuidDAr6zAMB6J420iwQ2EJO0911d+J04Jqa7MZ+KwGguMswENFU/BtT8gC
P3EeXZXGjI3Tx3vN+yjn+1rL6R9/YxavFiRo/btDyQC11b8oa8hRt7KrtuoGN75XLxeVx6DNK+Qz
WFeKzLAEl5Et2DQGkFOfDG77XFrDuBby9ePeGip+WnKmpXBTYWysNRdxXzuaxt/Ha3kTLmf1LD2X
Cco1OY22zKE4RkyXj2G2tLACy2SXraAELsyty6vQKlq1DOxqpOnXZ5Nss95fnh1hMAfhmQnTyO+I
QzJsY0kaIqHDuy/37I82Q7pAYMzSut1eBvaiyrXU56pgQ+XOPYE0Ogmv1gogZARL1YihOEpTPLa1
unNKzeRieScRYZCDhk2o9YyNsvau6oA6X280xQ/BDrNnLUAdV+eQ71P9j5BhMd+wt8ZTQjZQOSM5
kSQomxH/DER/XiUgCCmJLE/znv2M2tPwWcmhrLYPYOrTnGtdUOJhURkm0dyoz2g2bM2N7q/TNZ64
EK99zKGQ3sRjYFu7C2qUdmj1j3Jxb891g1W/rG1ZDC6UTIh6QdNzuAqNG0diSlE/nq8hlFM5sTh2
3BX6mMUUaeHUZF2WJOw7xR08Q+Ckq+CtpyiK0npv0qLnAWBlBQ9earlAStNkZnLSQ0f6CeGXbmu8
f3hcU69jFogytIaTiFQBOKuh/+0QPpSzUcPDfrYd2kjbpaIIS5WQaxxy5oYz72pYHIkWM4MLBtem
HMuD3Uw5DT2u+HoD5ot9PceKaKxsFOBUfh5mEUBI4EHw0wyU9XXaJWQUfN8kzbCL2RYyxRtlyK7w
HQtaiH4dXB37tU8e6lpapjxLvEKYMY4eFkmfcv16Eo/podocYpkqbpy1Gs1oiNhPGFzm11tVaaPq
fZAFmdizZ/Dqn/g962Y+2EDQj2j31w1+O1qMuCXQnUkPU29Df+wm1aRBpt83wTyuun+XR/XueywT
fZAotOLEag2GlKRBHsX+dt8zScymebearY0r7BOzTq8+DGqJPeEacenqs1b882oUv5F8/TqLrF8s
1v19Mm9LKwXkFnG4LAi1DBBlQ6fcitpLBAvprEDRcODBx4Bxs69eGnCnCjxM6oH1SLnzpoCUfhou
1x1nQIvWAY4pK9htCJmCErcX5nzQJvGLIz3cbJPsaYW9e8ZBzwC0lV0jRd8d2JczRneU7N3P64Le
L8gP+rvWPsgOHt9itzETj9wfp1lcW6ftXYBIizFcPmr8twqrhyx/1zL0kSBh4ILZHvQV3VrgGzVK
orPddOgxE4cokFNNRPnckOVDdpnJN3tZ5VdEvqunCsYs5jI+fWt2DN/4jdR2DYhxnf6dhYp1m5Vz
k7GwCUnIaiRwFO/fDv1LPsomWhvAvr980Gk44M/7ID5JAL/PrkMPILc7QNe9Yw6E8GNQ6tIQeUXr
tjEK+4sBHdx27aHIdzCGnQHZluyE7KJT1i4WuE8xKiYdhs5+AouMeHz6/3QDcIJziOkvh+CHbZ6z
k19QeQB1IqAL5LeYrxw0Jws7tUmTOUOZI2lSENXPK11W4HJ3TdlUBIQSMnnOrlCalUN9U56xbXgG
n4NrsoNBMzvcz0Wng6W757WGfKElkPSSLK7+xN0zNDeAVY3TNYDMHKUh6ckEmWEwHuZ8xVQTKPml
MxeLj0SOOuNl9bFPxbFQyVlEQMhafC6ESl9weFZ/yIw1KmAgzUKafWLZ/p88JEPBANS1P3Q+1blq
Sm0+Fhq4PFE4TBAp7fU5RSLzuB0msZw76oXVL0YOHwL98MhaE5tuGkUz0QmfixhyLyUgz7BMAOTe
V80CRwtsJ2Iog28y4gMdZDygwU5L+o4uJKIuUwKgTwVXDrm8jQl3A/j+k+x4xQS9QEAm4A/6hJWD
Wu+FJOJf5FcnyhmN+v+WjnWHAosPWcSig6YX/0LuRWlyWF3F0PHLUpPYujGguWaAlszOZBjrGnVy
IEciUIk9tZHJDrSblWyDoNEiw7OMd3YC0aYmXe67Z4JBhRnJIkOmtIos+WPF/7XAXnmRCjwc6aLx
Vey8anuP+tM44GZBuMgJhVR0Th77M7tAMq3dvMGdC0etEWMpTKOs2fr6qjQvMXnJVvtCcF/HvMf4
oWf91V7ph/xyf69HUmhD1DZxz3tCkuDVzr9qO5loeJrbRGGFTrnT6Sh9pK75Cw3J70r1orfPpyEW
M+XN7lyVUHnp1WJM64hd5T6rbikSO7xiA9KfwiUDf6fshd7WapS8rmXYtMgtyIZr+XdrhR1XjkU6
W45s3vkQr+utmz4fSn+prrqzC0GjsALLuDFjnTaVyJesYc++adxe5pZJ3eERCSUT0THiDoMf0kWW
QlJAo5QasjINmF+94gPC0bfpyDlJugbP6L3UaWq8DCBx+O2KZSjwmEyNKGa4Dg6PGo6hGX8OjvRx
WlT/8dOYYVUAOoPTY7O23vsG59k82DH5vrVI3ji47GWpEJ3e6QhtRg2Db16rrP6LQ91PCgtKvzIt
Q96QEMgF/mD13P/FCoU1l9ri0LaHcAvtwTHsjUA5LsskzehFFZPnSyryFvg/u6TkDbuDafoY3iQw
hDyYPrQ+uLf+G1rsnueEOaHvDW+NjtHu8z+iIUzWmxNJuGioUnQfjsMmH0SppZ8fSzalS8uDLyVe
XL8xfVIBvo2zBXIbhzn4Kk+tvElM4zJInfCzmS+ctxyd/ig0EQnv2/DVqfbg1fctEs8G7LzGPsSL
+CbOmvZ/3bDvUuRrK7jpQcalIaFUFKZdohH8i6po6S7Bf+0AaF8yzMaO9As7+CKN96AczjWES4Eo
KhcGPsdBsySnlx7AIVpcpijyYP8xsVbrbgzskQeGTMysBwpl8o6oC5gLEF8anfoLeWUJWkCuCtfX
1QlINrjOP1US/M3zs66+1g18M6DzsM1SacVQkmWbwas1B6rp97CXf3RseKRF5w83o3JQWLTlO/Ux
n7kPRKbDzPcuZXcgSnFjmc5Zmz0S57/x/1wyoXRJXF5Zt+4XO/X0XUIIJ4kgsZbHaV2CwsaKbLNu
xUp0Kmbt5/HU12t5+9mKEN0fS4At9NpewhYFWwzvUL/nwZL6VIGlgJLoMFxLJLs8N8YFUubUqMrB
+5wmnwiMiC84QaSBdWKIDHcUnnsrhIoG7Nw8nhQppksaADgWqYbhZWBKJdvgjfj1B6fL4s+aGFQi
F5+W4EVka2b2LxkErbz4p00mkCZx6+s8Sq9TyXACyzs6i8ZPZfTpeCEaaQJpDSgf/HXlutjbvHzL
TwhmyM/oErnnNJ3avEqR/PpSCuHg0CmWHsyQGdjKz2GiKJU5PYP5VUpurnY/GZui7xVaZ0RA3ZtH
eTiDxxmvU/4h6sRGYK9PX0yrW4+aPmpGldiTwfMxrq2jI6iGMz4nWFZHrNoLcsI8ExR/K7GjyNut
QxESuSGjxznLha56N2EYpGAcZ5WTMfAP9bYEDtSxz4qpwJei34HntS6dE9SQ0wC6yROVmTbBtUbV
PCsmLE/VT9Ce4CRTwcjkOyJZeFWBwvFoJFCi4hiq8bIO8PxPdz9KzzVQvWdv2vTLlo47weg20o7n
4QkqY8q3sojS5zVm0xNFQkhuxrKXjnwcp6ly0rjYjyOQjaEYFeKmjJWiwRgwCSju1doxgMTIkFBx
StGr6Yv7SRhhYzthL0B+Wz97orncQCpnnvlpcJVVU84nDg42yh34FSm2hSIVRaUP6P6ELZYeaQsc
GHHegj7NoQYqpcBir2Yafc/h2aBE4qSUz+XyKxdhVnyIzbw8BJpN5hUCopMUymBVeFOlgUASsMbr
OicMecjWMEcjVI/af5+/7w8jwV6LVVdA24QzlFvfGx9qzP1DRsMRKwoyfrq8mkTbR2t07bFqXUoQ
K7qfTtdBM3MJTsXftP0Cy+gbzxMWvUhwWD/gyUz+i6xt9i3jiVtH+APUtuQOpUUy8fzHyRWyMKnf
FOEQZCqkF3uFPlnmqK9PFgsfuWi/3f4tVuVqB8G97usNYz8vuEEysujrsVaMP2I+va3am+l93ZQH
XcQYPtFxXvHImTh/jO02QrVuqvZCTaaShu0Wz3Mxm8jd55qYEGyoq7ErOK9hIXiTpJQabTA45OlL
D5Fk+U+wg6O3y7oXjvk4atXm6tUaEWm274hdc46C+V8uWF+PzW/5Qh4Un3Y3BN0nLFEe569TA/Kn
8rbYGGnEJm4pAZk6ej5wk+OGVPZxCPWVi5uCWJ8zJubJpkE7DyWD3J41R3d53d2gnWjG2yQQKXxK
QQDI6jprLRW2U4eBG8Ivu/azIVell3kL+OPb0rt4LwXvC9AajogY4zzKl2hW6R04DosX3QtE76Dz
N6Z8b3BSzstHLiIWBQC9gJ3TTmjTNUr5JACsrI1KZzJzxz7zCjmd5VXpz+2JWgJGDvkfMn4YrLlc
Uct+irl11bVFP5UjQzzCHxEDggjCWM7+O0sg8V7Lsw7qFGT23HXkTHXxD9ciI2LlXba064+PwE7G
5YAfBngC9C+VxKlBDqtA2AvCbtyjTKiB83biHi+kieR4PbTrBoAbFgj0vTmCX8+bBYEOb2Q/z30c
C46OTkiRakGxpM+VQIdLUkdSzw5xbi41rNgmwMIq2KEN0RCN7eZBMg8QDRxVLE9WtX3Y6vvLdbfN
y8rCcJM+F3Gk+IL4UeXsY+SOH0GIKpS7XQsXjAAZeXHt7lYJq+xP2ACqoABJv6rq+DArZpgOu4/4
i0onVd6nSKOLH+sokDgPzPsLp1tgwD3Iz8LHVjG0qX24B8wsAvldEI7EqSGuHIlTeD3OaDlpA8Tc
g6HzTbjJOiBzAJ06mbUqWe4goDNd+9PxUYzwL3U7+F0fwUPZmMFnz1BuhWrwgjiDqobao+TTmYZQ
RcA++F/zbUKjGDrsxy8aaKN3CkP1dv22un2VnpsGtVJp+gfwPDNpZWfuegf+46CldfeabV5bkYVy
aUjCON1XogH0SPwVaUdgaVsj3IKxi2y9uOQj/HQ86NooUYIMwA20XARIkqANw9k+LhMel4SL2eHk
xRzmf63vTXGK4nouXnnnObQzJvvXYIO+HOjg0EcwJTvCom7zY9mjwA6Bw672557pPHdskQE6Ws5J
Gr9UfiFKlIbkulR8nJbS9ZKssXwUeUaiD3EoGV0PeevF5fjJdtNiOf3BjzU1J3MSsLJJVbhZbkr1
uMyggtIqCXzeEzSHKIFZFEpoyjJQ8nM5TzH2cdFm320xuh827UZkSuYTdiAsKaMP1BxAV28oWFG8
Mcw/Xnm9lfA99vGuPH/l7Y+mcmILdW8AUSw1YUkxxIQqt7ubJvyobLFjDrCkdj9VjzsmiDKesRs4
snDb6IgFZ9+DzcIk0uKgfr1uEc2uhu+c4Wwgow5bh76lPDydINY+FMbCpEQJEe8WnUlYD084YCxZ
ZxPHpXoZ8olExPVdhuhZ0MLi+IlsUtltoZpks9ovBOAE5HN8eX8ymwvvEyh8XWuy4aLZbSWPxEbQ
Yj10d7B65eZM4nTdjpkxPtO2WX+AXu2JpDE7YTKND1RqaPyFrdyg9PZWJs7xo0hqJphKnrwpBYoO
7i9m0SgYV8jTqmxobyFH0V2wPg2Jr5JV0KoLK2SNTjeHqe3v21HeBWDDacAjLjczO4PDrMeQaKm+
1pkkDHXJ73T9mA1IkUN9W7n0jYbE9rrtF2e6arYuXNnP24Rjzg+mnXtDk/vjbCh7yFCBhm0Z5+Qa
G8cSXxOFo5RqXCu6tT6RPO8F7wgErK7ZZqJ21C/4hSmfJwh8U/2FaK1lZGCqHESYWh4YmaYk9v4P
Xw3EpLKMlrz4DYH3cOjGVbSPWoXK3UlefruPVWzPmrYXvzGYtH2XnCQ1SAmJ0ETljaI0/wMMWEcH
+Lc5vD62Kk8AuGeGRcJKoyEpMcHLxQts2Ok+Bb+wE/cENmHXC5hPdnKoIHrwNjfC+Buf4i8z7RKO
iOevm4Dj1rYepaP7A7ODE3arqXZ9I98hBVzrJjLS9jlCms1Q8U+KseVj3oR6BsnDq6fShlWB5UJb
cIb4EgiW+XzOlcaDk2QC3iu+N/uNMW8RfW8NllhR2m5up6G1q8ewszKIuxxhzU91Z1q3YKh1ibmO
HjhDgVTpI7EesGrmAsxmJjV97eHBjRlpwNbO4na9UovOnDX8+OtMVsPiF7i0Stkyk4h1e2Pj7fYQ
sQPP1bf5c65SUzaKbR58/tjqyhOji0sSaxwFQsptJo4HDL3ItYP39S2xp7oLhhzq3jsw6G2bf2qz
5vzUCLBOAkTwk1cOXdIpR7I8DAJ2mbwIAQ4FnOmXIfjmJFLx6i+RJWMro+3uschIqCHBRIpipjjE
hF6ePbGC3jw1hAgOU71w9owbK7QSkJSB738GufNXgFwnoNX9UHdraTyfyhb9WGyUn/buSFRzSRt2
54lPUjaFMr2to9pmEAjIOIDCzQ7Pgq0p8mCqD+rw+9w7n7doAKdTeuitnJolNNthPHuy8+i5ju+V
VK0fqpSA69g52AiEiRJc8tOc1g/nthwBKA9xSSuiu+lTd79dQKiyvWIwddKE83IWhQhlNGhYaKnd
2GUrUviTtOki6WBKdtZpXvNuGFFIxISnORd93XDReCFMeJ2u61BUDdpAeQt5HbeV16cCb87VVYMj
FwNWs0cGGBXLDEJudLFfdleEuFwhyjldx5XtimeRCiHnfo7eSvVweTg0irbiBKaOP5SQxMYiJRJe
rkTsr5XfK1vMd5E70ccxZIAvB70Vh3gbRiRUfNP5gFDCTkAxuw89m/HICMDgZKLdpySev1fSf0GG
XWf3KWKRy54RHDLxJFJfl2JgTJ+ysT9xeJkD0hD9Sxuh6HIr0nKPKhuesD7zYtKZQ8z9Zn7YDYB2
TmMbrUCIvcigqy5W1Db7KquhXJ5g04jy1GGDcOUqSAv3L6SOxOaG4e/70FwAAfek53/oRlqmzTcV
1pwbDI9C5imdWOJdbup6i0LHmmRmzBuWO3deohKq9etuGXJ9ukckFdffi+zzAgw5slNeWERzNRU2
3Jg4YvGSF/oDSornJNVDj8+Cg3iuHYW7ktDsZw0r7Fr74Inee/XYf4bSgQ2dyxp2QyL5kMMYhb2a
VazPUUQPgZfgu07/2hrvF+JO4y+mt1YAjlx0yd9iKfCP5ihGPbeB055odhPIo3zKlqkkeSquS0To
bC2L4ytE7txT0aR5Xxkfs4sb96tHn/Mf3/1rYx1lVVS4fh0j8AKIbazfFvUdHvqNIigLNzzqBjbr
EmWw95rDnqaw/wCOx7WPGQN7y/7knEfpUDz4dqE8u278CPM36kx2fD9sayJBzZWtJ3VBQSzr1mWZ
CLjhxqIeqtLFFyBRunTLZyIvZn98w6HD+ASjgPqH1CdRejcWDgvHwEm4ZaHxgrGnOE4Ky3M4gr69
66q7M6toOJ6NsVbvAPbb/srerSw2I/HvNCyGdA+POzD4RbsSMD2cGxawEyb/GMnMFwBNbZMijd0R
JtiYG4yvDZXRq8Jmk4T6sBq0K5JonyueGI7MeA+E9h/wUxwcGiQmKLo3rCXjlVZCy0YjEmM7Yn7Y
iRpcFFRfo8NdRLn/AXe7K/53iro4uBYG4JiHqRGkglLTR5R4CeA44QmdPiaE/Poa6sQTyUr+J0FH
hs7ZDeXq/Eo7BQojodhRJS+U0YE78p/2fPdacAbDCtFLzQ17mwc2XwVQfX4RMWlTeL0HX9veWxUl
c+3SVh/ECU2aFvuGVIj+9ywQnyyAOLIfZ1yBiNO9p4Sr4ZVfxX3IULcvCa6PJA96820JP2g8GeAT
q2HSsDtnfuRZK3L4woN86r5VG2Ob3ZFprq/WgRt5WgHd+JEdvC0Fqwh4jSYoZdrzqJS/8P+xexyP
vco2RL1QcTgz/dhkoaVVv95LurfZACXaNCfgbyrIfXGvTRBtr5nXk/jGjUqzfjBb/0kplWQX87Ur
MCA3oxdytvfh06pm6AKH8rkwGhTTqp58QmOpq06jb2XvVHqMV3DvnT1JWjIsIQnqDvXXn/HKQ7kN
eWrJppYFLnOtvXsiTwBbeLtEH7PMLY2lMLbGNz9Me+2jKInxP0pYEugq4qnk7ZmsJhXbYX1Cv6yd
KcNir0LtiqKkReuuQRbFxuSOWJV1Tw86XVVLpAOSeRePoP0M3TFUSviK397oJ2EXHb5kdzsjqBmP
9l7u0iWlDFTtq673LQL8m+rSeAGaaznH40Ot1PR2hYBbw633wRwXdq2cXhy4A0BvR0l5jfmoOYS5
c+Uk+eFhUkrTQdUvG8wruH34uYEWP/DxOQbYksFgkiHpZ1JUrePl0eXTqvHZXpEHbisjz39wW8EW
GKBn+Lb7xEOv6rFVuyYhovsCVjCQzpZi0ZdfFoWZhtdg6sKKKcqHw19EaPWPE0t2JxRjXbZXdQ4P
cggxkrfSr9uMseNf329wI4OcKMpItGeNxWn/IlYB/jrDAmt6lQUuvjP0Ao/KcHwpxT6JJ/NAJALY
tfQUkQKu4qI50SRrAjySomRvoCLsjwHik2RTnzH039O7BxEXScIiXIwDj4YEr2q3dPAidCAt9hCs
LMZK0BNdUzX3Pr6xAItGngHrldzUbAYv6CLI4T5AC6U/cpFyfjsefMwkl65Ozc3a4pjlTvtTda7s
IVvbb9uw0gPfSvYLsD8qtHTHMGDSfqRlK5k8LSgZCH8xrxKfv4EQ7z+vgG7NtzkjdhuVUHrTckDH
acgVmQk5qiw5+v6cfaOjbcefeJ3rPIWQ+bUcqubiYiimKyUxLZqovegH645g8u3dI4GobzfHARSM
mBPsusfYXtE3/iZXgYqPVO4Ih/6opfM3KlCDZQ6deFgASrCzu2iVPKod1TpKpDk8wqPY7n6BQhJL
+i/yJA2pd2wfAo0qXa8vRFVsluwmJf/iBMGiJHtA6u3RbzF4fRx4N7aKwUC07YxzXnfBrOo64P6J
VNq1HRESq+fQYFQ3R8HI3n4zIBD5kTMat9eAVAWCx6Z5iwxkI9dnkp8vIfNZsQYk2350dryVZ7RL
KvFTFe6fNDkrrK+qLWcnBoF5iR9lzXP9Lj1DP4r47DhG1Pj6MOOX2nbkSkndHn9cQ8n2Eaz79re2
IzTpgBT0yoTgYUnibJ2mipGAHz34ZV8iqIKgx6P57xmeKrv3NW9h3sF5ZzZrVKjnBhYCT3hiINdQ
ixwSim7CYJAx61UmpXpyKaFRmQMIZcAtIDPZvr+5C36rhdYhsrryZC0yh+oqGy4O6lDuINVZFW22
4KUBKdbaUifFa2Tn4IgzR7eyf2mAiwuOFQ9d1fwCBShtbvgJVRL+PbkCaVCgpiTNBei3RSQomAwS
j+KRMjoUri3Y2ShCvkiexaDz+1XT3WDWuUqOZoAeteFqU7TQpQozBlq6xGNzHwkMC39hU2fXNs5n
k123H9s7dF2/RCNoPfvvMjyenktylz3SkRt00bPXPTxM2Omkn2r7EBK5ecfJJANh2+arwEA14nE2
bzWqZyZkuFgHc/a4gtGpOUJEzkVQjsJ8kx/I8H5wbwWMI7IxAugEMzWjawU/CRkPkyk+ca51f/yT
9+QWjeKNg3HZyCiST5B87UHcI5YvFAb9Vv83xMQdvDOCfmul1B3gvM9ulxQWAyNj/gHYrhAkaRxR
TLQcrgq1Q+9UoG97nuq8yEevPAgfSFSt5/jm0J6n5S7cCRVGQ7UFcva5HAnZlSX5lyZdYIX9fExh
2VPCdlUdAY+n9eKYwu9mUSpPZJU/+fbpqmz8UDwv4D8KdqjgUI5BH93wHXgv6SljhMJ6rqknVRia
RaCW4jC9R1etd11MpbiDLWnKrEOUaaWr5PSy6NDWFetTsoqtxnJk/yazLfYMDgMyzwRr6n4ZkOb/
nB+3MflvIyuSBhVO2ymgUmzR9UEQdjVlG8liU2dYcVORwQhqHLFTGt395KKKVbvzf+BxoyXOAizU
TGHbDI9o9pD8WpH0pEpP6DDRZ+gd3x+OUPl46AdEPAvdvp/y5Q0QBEMY/zUcnN32ldi0jPVZuX8A
2fMz8kgUtgkWdTC5+l0Gq2IjpOqFF0J55EWxIdB50P9ud8EDzhSFQjtE+p4+4xXzD+m0IVld5FW9
QvILtLzooU45DrHdDPfmWMb+GsiB28RjCRtYUuAtp1rMXNiMelMLfPmsA61tktCJO467AcrbnuDJ
ZmWjX6bNH6ghf8uNxEbCbVm2aAYO2ADvxgGyGZ7YgPar6FlhPgUpiuSUzcMVJyaahaO1sthyFOWT
TivHaI5D5AYHZstYjVbNmHnEc8YhHusNkIYzX79cT4Wl7CuOH4q4NrKugH/QiCwVc2wTz5hKu+nA
Hq2tu3Tl0ef6AWSN7TLGA5RIJ543O/h0WXj2gficd0G2E1hIcpU6sxxDMAw7C2JfnHF6ZPG0S2e1
KWrUShAZ/61hWTcoSm0czEkxUg1Nj756TOWYZ+D6S+laHl6KKHmFcJxiOJu7cEenV4KIN3ls5fvN
T+zSH8H7ZJLa2sHMJ9M7X7gnr5RXwQvmaynnDL/6W3uLtgRRECSXpBikZhRLG0R5fnUbMrfS4Jag
Wv9S3ydy8094HuC/G8ubaoi30mH8qpR3W3qnDXM1L5lAPjr8aRori1I1M9cZYDKnwRXv93HZDnzz
TmebFHkHkQU0iNDQqU0vzvgbNwf1QdQf02pWg2UkKAwkZ28sXaIbXR4RG29dv4FQGB4vQgThjt73
+klre2SKR+3T9wBmFA3XnwhKoTDY9zwSgaUYCbV+wlqKEaT9NKy+L24clzQXnzxRvx1Q/E6LhjMn
M1E6Bd2eD4K2NOO5PTT+4MHHdY1EeL268gwmDU+15Nh3NtPhgp2pV7w2igqcw05gxZpIxgM1Fxes
BmQU2HxeC4uLUoeYexXsRkbkcUzmeA4aT1rjYxELChBLP8d5xCxWxZhhkQ5dh/gAugh3clYMG5G2
ri9bh1ZNctAxWkgyJYH1Yzjqyv63dsdEAzMoR8xiWQmkRA56Zb4GP5XXVGYr0ERfqFPh30ahJwBN
TZHERwn80Sz9nVbGq/6KXgQn3uM9/qfOztX0q5CfP0qiTTT65oqeRQjheZYCtYpe/zC67TJ0Nhg+
bEWUty/AsKgEnZbTjVBgab3OMWKNNZN1nxqMlu/GEo7NTS/XeO/z3tbS5Io+tkyPXkwOMdNxa+RN
TjNLJHJS45oIWhXb5FWhU03klwNcLoIBZRcNRljTmfDgcpX5uiEmJDt0WHjb3AZZ7solWNHvq3F5
K+Q5hIecs+lIjSJmz+kGzIVR5YjvEH9q6GLEaYDwYMNAarsEU2vMcxifMugkbb/Q3phYvvsQ5O/T
7hEItFQzQ3RR6UtUvoQlW573MjtscWHcrUYBqa6QpDKPzQEeZTSvGSN2QOukcWyd1CXLM31/3a9l
YBiwQpA62QNnnuVD1wV4WyU2Cf5hkI2giM82NBc6ktj6g1LNDHzYUzk9IjVBzOM4TuRAnSQbWd99
G/Awas3h5gI9eIBj2E0WaRAcRnKK2dscfz9bQONlmozP55cflkZPuX7RSQMH+TNWbKWicUbHdHUw
lOhJUe+j8cn4hhs5xMnaVoXphHXzZNFil+PhnYlIQxxhnj91luDPue4ZqWWj02f5nS9vhzGoVCxM
LXiZpF4hDhNxoaYnafwK8DSr0p4m4x6qzguyBURv6wMHcB+mjrFJQWdPPDKUqKX7yVZYcIJgXrhS
NuE2AbhNSGPN8L6nL5VYHgh2U76ANdVbUXw34UEvS47g8+2DVan4rGj3C+AibIRGkcVvP7xuef+Y
6RfgIKWcegaIdjGQPbwUTakfDflwvqQBTNZC+UUwCiPkEAMv4/aW3ZNkqKHLq3qsCGcyc73No9nr
sBFXo/vJhpg7t8wS1xIdDKbrArd++6n53+VdZOc8/rgM8kSkq4x4IMHxUoNkrR/jydqyn5slMt5E
tSSSCZvy2VWGJPkl1BOn502F76/UaEzuzlEyY5xfxup94mEcM+dODKVz2HC/q4FRqQRi1kFXjgz0
x9Xl8OyjIOJ9YN7Rn5vOJSVFa61nM3h4ssqillLO/694g8J5rQoWG5QVZ/BcbtZc5Tf4hjprkZDV
0v56QKJOmi9YeVmZuBElGrBkD+BYDHH1X6LPzo5EayV2urqGMYML7/ksyNvOqd4fkhgRaqt/I1WY
rulxEH/svxwskWopdxiVji2odasW8b2k1vCV9OaeCSgXRJThvnpePv7K8KmgQJbREvmDMDuUGYKa
j+dVdK9S3kvkzzBB0Z0Wr/utlw+mRH3/99I/CWNao/+Z0cI5oDp4ukclWm0b2B7aFdcgzNV/g1oF
ROIy+SWlA/caoqk0dQdJlBvWmLWc9tRna4Bij36bX3Ze5QhhN3j2h4E6GzFmlR6HCg1yqu+5Shmy
0lysEBBSELP9+wx9Xp9yCcfdD7Qh1hpxkGyF6N6dRMSrlxeHWvmFKcG9StyQm6SsFiGUVWLUarZD
eNkQa96yo0FgrgLZ1GaQpT5XFkxeuvkT+smlHfN8uMdCRhoVsCsIFURfPp+ELrZKi2mEhy6pT2GH
unl8yeTfuHS048lSrcI7NSO0wLrTyAB598fIlpbETjbm9G7E4HaevTK8wZPrO1rVct78GFFrC3X3
DIh7anI9aNeYgsyINRXhCwVHbxrcJiyqaTpmasqq/e9szrRdvsAHmKzHNrfs1dUG2MmusO1y5mXp
hdLCg/bfqpIeE7V+FCOk39x/8oDUPIXkh3ihHjGmTmSA29dRY27W19TNBGpZEbO56BzaVn+pG6o1
hJ74qjt3HBD08jJooGN3oEhIvAOgmJKlGplyoO5cxdGXjh9o8/8FaYQaNaPvL8ETrZRDwND/SGp1
O+8F3FMxUqwwu23PRKYcqMgWjGftdNYXs8b2jqXuFbXVctJyooNEnz/bh6pTZimOyLUq78Ze1Pwp
YVfz7w+mlX9bxSW1fFuF6b9Gi115ZDVxIksDdKJ684FOD6ReytGXw6+keNxOY60J+52wu1MntStV
zHjeulcPMaI6AHXvYZe23VLJjTX/bwf2grM3Np6tt0xvIktWwZYwh4umqrChiMjYAF6JLs3TOmVt
vDDyuJRP5RsG2vYMj92g8AyHHCawD4N7ecadsRTkqupx/RZvG/o+SR6KbXZxMdwwcIIE8sxmcOsJ
5hSmP/oHi7YvvOb4BDuOOnogGgpZ48ZsQ85dFw16NnpkO1+n2oD3dkshmCj8GnwhGtHcovqepScK
1nQNzw3mqs1ITi9QN63zNQCCK6577lx8un7V8yOPw+Wn14nauj/ugLxdJAAbeGYX9bPd0MpvN6yy
2MJpZakn2EOI5T1gJdFROya7h5Nr7dlNQZFiKKhmb+lvMDRQd5RogRHPJ1rzrBXIEGgYfIHjeREv
ogLac7FcPRv2J7YvA4pY0IWyWWm0GGlYukNctP9AkbaYzLc0t80povpiW9lzP01KoJFruM1asMaP
8xA2cmz/fIcPGZrzORiKWOI8m8scGoCaC/J8ij+zUcvX+HdusvUWiniDQVtKjLFpqpb8ES2KB8PR
ByykGfdEwIUfgwkCBEeSgBrGeBkmQ4OmPXApILCDwy0XcVVfHrVVoujdkW6fwNuJsfxeXG0axca0
VC0gCv44zksKHRk61wvA7emrv/y26JC7yKLqtfV++wcNqPQxkJBxDh4ZMWj1h+GoHPT8uzQz8MEu
aWtz1NnawKRKyANctKJIFDrgPqaAdQvNqE2nwR3gIpFimtHkxK75Veu+sCvf8xvg4dCU5ZiDED5p
kleXH4ZqoL5eM/TAkgGRgWQv9ZE4+RVfR68pibb7RsNtZeKfgUKITmKef1IWMZMcmsY2FH6QXV4K
pZIFroQP6p6+f4rHpfBfiJYD4QWFMJ5VDZbUJ/5wXs/epgy0Q7s8IZvXYecmRZcm1ROYr+PHA/g4
uLbnds1twCzdXiArn8NrVkErPgawRjDUyy5S84DUiOYqq67w2M5MxI3oD1hBx6wfKpcu9XXFpAcd
imzmRU0kO/Afa5iWKWt1+1zlWL6B2CxWJvhXrcNFSANixyKqDtcbs3u7wXvZ2r5vs6W7qJu0fahE
N24pN/rhBZj7809twzaCQQ7QdQwtt7U+jqRcZAUpMwTHzQt8pNKXVGgF0foKPjtkNouJt4eQVTAb
vHG6jpurhieSAd4bK4GvV0KSCIVKl8mmneU+cLoSXh/IZHG0NxT99Y00hGQhPLIBifi4eMgNtppf
HDrR8I1IWd704sPDtV2OHm6Bu6AM7e1/MqfI/RGIzGMrfAfEVDOBFLOantuk55rAui0/DmSU6YkG
qEm2Cw6rn5IwNoaTOuPeIL49rt4559GqukKsmoENcRUTCxNtCBwTV/BdbwbcJx+j/VBIZMQkqwev
ZJMttV6x+MzZ4Wc0pfbJ8im84kkAaFUdj8zTtGso6S+vwz5255U35NLfkBjONn6FDZjbqcRY4gvg
YEX0Eoynf9YcaoSSWwNqxaGeII09cUweIUiFeRqV0HA/ohGWt8Vi+9/j3+YsVLdZG1DsE2hE7Jru
15wgjPSaClpf9sYvQQwzfRUHcXHeYM3mEG/ajQm7V5k0XNsmye9iaovjhd2Aj17Ssk68e6Are4I8
9c4JIdWG0DAPG3A+nqfAmNgfkD4lm2c+2UU4kHO1pv+jw6rQQHhPLiVG8Gyz42qRW8e0ikUsuWLU
qqWmD39+x98M3QfFZdg0e46V9TxOXXffPSVO/nG4L7JrRvbt0g6rxyxTK1hLpH1w2sOEaC0M96Gg
g/SoHL3HWs+rXoEsvnX7h85q4YOM4wCq+P0JIyK4TTiAMLN8OO2xT/xpRkOEavJTJxLJBZCbcIgt
s0O1xrwionI9DtrVc+4uQC1aOh1/gy4RhP3pRf729qIoWViqQSABVNufXIvI8qvqt6+BOht18d7Y
+am1Xeu7rdEGG63asQWkRbN0WJDDsH8inaiFxI2pnmmAwF3QfSqcGdAAqvyFnm4jp6uVr051W6OP
hae6uJF+xQPJaNGVXbSSzQObUrEwma5aMnaYb/+f9DDHtCRlU6O2bHk+yz6KW6P/diOUFAa8QYgs
uht2VA/OSVahCYAZDkEHcYKvpq0wwazdx+ftwTYR4aZRzj+YnpxxjA+M0dOgTgwZEWuF2tXZegyN
WbN6sSbw3fuotaYpWNDlk7bGCUnFf/PCqVnZ72q1Ld8bdXVlhUofCnjaECDE91l7OHRwe5RFxZVJ
3HN5/9JaFxb4UEgIK52z9GvAiEn6ynhr1Z5T+rkVidtVwC3DNID7TcLLPLPQ0XbtrZiL2jimfm+g
eQ13vrkaVJPNVwTqgDQnSNgGKDD3w1eQDU4nuuASECSygq99cpioUtVdTUmr8Dxveqi4nEwYRHtI
i0c8BxM+sP1QGw11hZ9e9i0zbH8w6WGpZVQQgD+nA5XrG1LO5EuEq5XhW9e42bSYkr5u7DgznSY0
zcp0ewF1c6vkTWqb1pmUer8TgMZ5CR5l+ncNxD2d4tQz7NzK/1ffT8a1rFmQgxcdYj4ET6jj5WZE
rwIJund84+y/3cxZM7p6sGlO9XdgURw3h+1ZUbUfa5aUdbKMmG/ZiISRDXsxX6H00gqDKaFl+S5M
Zrf8RgD7Oyv8vTC8v/SRKrkIGvjwH5khWcBXAi25/ZsV4jrgHyhUCD+/rslTXeNfKOcOJUjTAU7S
n8DEOHQcpwEu8ev68SkoZ1TNMN1527nZy1t9JQsKMJyfLjw0ZtIst8sjVAd7+cPOJRjNqsWLnceJ
vR8s/72pVcAHJqJilOtlEoKpnTHOhSL3mb1nega9wkJi/D5lm5O0rnWcUwKxJWTHPzb2stLyqrDn
PqdvKXnzYj/KHv3gafeYqTu/oW9js8N46lGycva6dKOfGQVirOg+jPniTKSoES/uRXCsdwyYA029
OwYE0KAAVwk+sd+wNdfOveNnu1XcE/RKo08h7itt+VFW5VQrGod+mLz6kHLyOw2inqLO1rKgPlog
RPDgz14/9jCOtb0Y7JkiTd7a+L9zTwHZEZ2O47Fhlf+PfnWd7YUI1XV+EFpWAKxBEHtDPBu03BQm
vOpsjTsD3kErRf/nu6d2EAnwQ4jDFHXsrynL5Az89az2c8iK6e3tl4uTEyYkpnoHtxw7+XSoRCED
P2ELWXm6rxdTmlYgl3H/PGxpdCW8y86jwt6/TrL3bpVMg/+AlCtaGRcwhgK63AOmNkC0O76dO3+y
yVact7vKld0cZIXa2xi8m/txXMSmFFOvrxKMveDlE01rscu+RnSDmhMwF5G/6gGpikVKgXiZ0+Ne
igDOskP451vecvluVpMVvS0z+6/d6V0SEg2U9oYtzwu731QmmvS/eXf432KwXSCzJ0hYDl8o6IZD
TOblsrRokdVtR7xm67JdcdMb2er1LuHTSL+htFFte10hXWrS514nqqjtVMMpzWywOXogQxwz4G68
HqosMFrDpHcpBly8k69dSPaWChRXzcsnksLqVaFdWXsq76d/kWLHtl64MHLEO8bZNNrMyp7YDUJH
Hylkvwbu0cAWiQTP1XwA9WbUj07rDBUPLXYZOShKSpIUG8Lf0wfpCRr8sVQQjVaqKh8QO9G8q6TL
nVfs0vTerWLryMo9vNLqA6oWIujBfVLtHJGhXDY7VNi6okYRSPjhnIqby7Z59BVggtq7G/UFJ6KU
MGcVJSfOFqkLzssFbsSyUA/QZgeVNrpeer6N3GR1uRvv80cN9XTe++d98LSEt1uu8CKra7L0XeV+
gicu9J4Z9Iuq8L8gY5MFzPfH5+Z/gAHDPCc3OqwGUGkw/12ksBTHnjuYVkwTLPXDATcbpuwrCyTd
dlkvKO0eZv/4QIJVimmh9fLM7DIyrhFz3LLanRNhS/vyWbBWyCAIj7QykOCs5h0At1uKsMvzv31m
ptNxAAnwE90IZ2TxYz7Dwh+Zg/mCcNoSUe2aaAi+yJsTiyzfHjek7XukC8JPyyFhkn0OGUTHHlqX
qocdzY9gxnpUD9yZZTEbhblgUeY8eqezkzhKbFqw9EvPf+jN1XFOV2Gd8ZUjGqqtBgQue47K5yMS
a3xevm25er15jycLZLPoXOSYYZALOlyapufEaAO2PYUxpS1TujQbLs7z2OlJlNsEcV/u6FyT3jjJ
QclgYG+Qv5gpOkw2DKIFvfiRmBFL0Klp1w08V2HtpJBx//dLiS/11gpiu6IBf1dQvqXdjvbOsv26
BRnQ7knTI+jGVzoIic1J+wEaTeomSW2SvjkGFQUnB+1SmfYSmjYpTVeWAM4JAW9mbG32N+cSQywm
iRFdli2NL6gPESfQ9ucsQdAGrc2+C8H092ys6mwT6162cupZm99ETIja5IM9vLCyhrxXru1j8zPh
8f0lXE4SU3XijdumSTcVnI2KutsgdJ6F5l9OgbxBB23x+05Eu63U/A82Jl3ScFfzlt2rn3H4fwdV
d+sYjoGHFCNo5AFcVHmVHhFkq+OWJgc6z4oKxFJwKQA9urF1nhXoHbTrfdEEh3ZVCVNqWnS+eC6/
G+DiokI9YY4Q8uR9i3Ej862ekALrBvJQl66UkIaLiIl0piUg4/X6RmEvrlpIV9EaQBoCVRQzaJAu
TwE1lhxvMVm2uDAFll6kuNBeqwGM+HxhoPywO8e2ZtViKInH6gjnT3C2uT4KU5wZgvt6W3vsRSUy
naboRfRZyMQnOxWQ/bbAsLKTnsCy02loML1x78KyhjqAISRAEPjIA6pJy4+0/2fY2VOzSVAX0Ml6
Buj/0n1qHkzSSb4vbswiwsBp8zEJK/hzB9Yt2h9EBfzL+HSP/ofayLrkMN6brNEgD/AwKOzL5Yl1
StTHhTMSR2606qyoo+RthN2PKPcbt5MRELZg16cdJ6MnIrVPHrjmkd/ImirRQfc/0hCMgjdd7X8m
yF9oQiExOwoM1cEZgjPNmZ0pzEMyYhIsak5BVVfN+A/NCgFDJNwiXPl5vCYMzbD85VCxirN0FY/P
QqhCqGsc/SU9h1dZFsUyK2ByhVfWutKCF73D+3eebDau3gTyvtZnZK81hIRCtbtU7tcl0FsUfSyf
V8ItVm13T51UIj9skl91Q8lPFyX2w9GQNdPW7a+qQ0mzihHax/rOROoewWgsYMCK6qSJwZPwKTyB
r6zYsMxeSEy6OljpU1gAlgDME9gwxwH4GGUw9sdCXaRqfK0uCjpkkE2bdqVVOptKbZplwDFDxZ8O
qQk8AuvvYAKsKXdVOm/U14YKr610Z4H06QsIdQ4CPj2y5j4iImC3fv7ZCFAoXQxDIGKu+fGxSYzM
ZLnltR5tOaKut4YjytXnJKramtwkln/ldq7MweF/8F7DuF8Ir1uSS3TcQfLg/4fCaJaap6jEh9BH
dI2WYwtOXaO0OiMoWgyDDR16evcLvw/bSaf8WKD4OhkuhQLxxtj9qtm26OVGF9eHDTXTNGGB16ku
ERhM1ESzOtWfg/b44bK3iLDioSMF9vBB9ygDzG19DJ7JH6q+2LucUbAgMFCTR2XKkVh84I1sKx+E
YUQuiw/gm3ucDaJci82CajpvWS6x6HGBkbXYyQxXrIF3/Ee0FU3LooUmuhdhMS9XOU7RfI4MK/+f
EpilK3votXRScZZdAl8SiQmBz/AUaEEwcsF0kq3uXbd8G8OBoFmKLFqhMiiHnLmbqbh1RoyosVSA
wtCEXYMT/oshMBnxBf74g07wv63rtQATHrTxXc/hKSdNIQzqjHELIee2Ztq4T+dnkdqgoXtimFDR
YCAWelW8VH0+fx5IeBqnKM7fslK/vV8rUYFsv4sutZQt1SFdmz/rWE2ydEzb2WPTr9AUXd1zDmyZ
Po9josrIQpExza6b8Wii6V+WWtQSgzB66FaL3lwS+xAaFnBdnP9i9WfOtKBG/FQKYh/qtJkM+dOz
qSlkiPG7/cGk0jrhffSdWr/+GIdqNMgYBDZdlfbzY4gNTUhTehFfkOn5/+8I+BzJQ0540piKTPrE
ndGet3+iCBQMXbt/j22h9bahZklHfsXNLB2op4XDnGmHsz27FA3+GfFoZyNVWQmGAST1/h2sISzd
3s9jdb2BhCII5zTAiEpzuZyXHdbJNuKm3NXjF5H0HYqJSVEU70N3RbqwDcLdEMkOe72Q2yjpeCo5
QiI3aeE1JCP8XsTLbHC+BLVtvWcszTeBkvU7H+C1BBF1zSeg8pLZ1+zJKgNh8SqOE16UmkFCzS0m
bG/qiYHPCLwWYboSJIcKbIPDB1T3xtQWO7+YguvVqzutqcqFb7I4X2tVzLuo2mcOynZnNN7ry92X
jxqk/siXdit43l4JEweQxzzmYRtRhaiZ9icFKMW4t8KQSDHOpU8nKjPa/UwN+XElO4sm4ERRXgud
cwEmC4JLeLJzSA8qafRbzZBv46ZNIzTkocYJ0z8YCGtjOAzLaImSZyy72z5v1+9+q//iD/LzmWCX
+spHbB63FCiRziNyHb2BAKg9Xo6k4/mEH29tGGFr2KtMfuIzM7JizWtPut5CcM4I2/qQhW0DtyXI
FhDWOjMJobFYDULKAYmAQePLFzKFchgQaypCQDWAOhjEDo0qUoAO5ULBCzq4uCVgwntW1dFVDKMr
IL/njMoFc0A80yDbC/rJDy1FTu1gLNklE7zkiLP4eWlwU0+PR2JEEctAcNJtw5OAoJ5vM6dCxnAs
BWhhYnt36ru18vVWIQOn4pL+9D5ZlkuCZp0ZeTuATNhmfovseR/mket9z+WbeLJz7dCfMC7l/mjM
LsUOAwaX2Ykb9Yqsww2N1L4phtS4I7o3EY4PUtnhlyJ7XNbjANECzSRz0QcI4/8JQ+UHDw2Akh7M
evy/Ick7cDdfOLUYX4l8pZf/zJbj7bd2SDhCraspuKnaX16YeF/lyZb7Hnhd/Am27SkF92Xerpt/
KiuI4fcp/LpKMp9NcbYyo/d47iCgrdqj7SpV+MmIdEWMN+yCgc5UyckvzBgLUOkBHda0rPSUiMC0
VScHid1zrKfEj2r03l4OfXv5yvj+3rBKhGwvqAqRwiKGLqiBG9Ny/KtPnwu8VOcwC/3UYxAmYily
toEg55gMkLHClEWHE/XDP1zVKyaPli7hu8shTzGamOtDxsaCg++OeHoSE/AOHnvPn/iCwQn5WUJj
TqaIqE2BEqV/HKpQoUJoOMRKkaNrNDMX+dNayC7FRvflXXiIUAjDb7+ljNy4Q/fgNDuXb2yUbo4P
ooN5HIMY6FwmkObE/k5sI9TthReZnbgtHuxc4H2Ao5tqaNfPZwIk3Bhl4jPN+MaK4AUO8aFnamCR
GhyMoKxjfG3uQ6VWZOOKSgiCiWPxDmUm7zkrO04EqCraCfBaDwSWD06Z/+Z5a1+yUvpz6K8XYoyp
NcMlHy0we2WSPCWnKSobs1YdGdbyNPx2m/TSQhy+a8/LT8kxc1cMTIIGeW4MPHcbg0tnjoyaoLQx
prOIj1s83mFUbKvBqPfrIBje8wn9PDeVwCMIXGvEg0B6xbLk+L2LDjiDfV2GOSIsgwEB2vL0alkL
o0l/OSTdGfO8pG0NVzhMLj6Wf8DEHeGgHAK/xtcKpTU6Gp+8SP2oUeUuI+ThvRm5Ex/oUzhVRgNn
72t91ohyGsTAo04k4KyKaA+gQ8QUS6C+cgHpVSrhWiGnIPtbEspr5hOoQx4DBDk7DIcYcFDQSWuu
yqpr8RKjF4dRDSawoD899sYcCL97sEEH/wvOoMB5vAATlCLF8oW2tdlGR2KuUJvJcf3ZJMVOqzuN
+uAcFWtRWHjgqatA9x5Oop0c6u91YAp3IMjK9zeykq5bD5ayJPyeUl22MhejWt+1zvP1KCkJMdP+
2vOLHgNKSwoXo7tJLe2igLD+5tDo/gmRUmMpJ+cSyYZlCH5rem3wW2kz2s/pFqRdL1hTIEfixSQV
UkBna5eOpVBz2vEemu/KzcTzHgUgqyb9+d0KyXcfAy6v8DHVdLFOCfBDyTvyCJR9PMnzwjki5HD2
Qu5RR/30bC+uX+PCVQaP0m8cq58uObRc1BbceQwnzR/cQoIq9mrakjJNhy9fahxiNs77nuv3vp2Y
MC6ZpCjjlPFnn+kvXfr07nV8zaA4mz4cgjGaYyXt4F/W09vnCgoaQLsvAQ1drsAIwlD34jQH4Yb9
VE5gsq8CYCRIVR6G55mONjPLlz0OdTJfl7LfMvyg4CvJlpxEsE9o4dYMl9OI83phmA0CMwA/7WKL
R9ldDsPwspPQw7rQzESMK/0BOF2aIPlvplGSHTTeRCl0wp2X+rtUfc5B0oK05Xl3gYz9fi1o+GSM
yZ4IFtOFoYttk2bbB2cGdzXhAY7C95T578bVOkpCpfLJxPnq+jKNfMjEbwq9uA7lpiHBj1iSVjYL
5NHkMy1CazRHXsm6izMnlQcRO2XH3lUwy8v3svKehojDBXJxNuggaG4YKY2cYVLAfdT0YQolh8Jf
CMO+38glHLHvKtLepziMiRKbi2h935Mdm9D2v1x0tHOCoBKCfoBpMhCDs+L/0+qhjCxx8yLigmrC
77Zt97Nm2tIVp/WRjsoJzIVu4L/I4nIOKdF0dAIC7JA5FD0Y0pA2br2B5PKa5WvdmMsCWxplGicu
JfmpEU8KbTsumSuvKYVSrn8O70F35YuCWD2siEWPw+qT5CLkMSNWiTr40hqsc8Q9BzuSjhMRyxpf
zrEaFSDXVdPlK+oKJkFrBpQGR+KGLSJhnMeH6Froe7j8a5nSNVZPksMZv2UWSVajowfrVOOQNXIr
c1gfvg9JdiifnqSC4VHFfe1b3YXoVkYI+qnMC1j0ouuGCdR3c1BGWsQRLDismoOqoq01/NDdN3E5
0dF8pLfr/E3HPflTz3PsYz2xs4uO2q6a0f+v7tjMWepcalJxoKHkbK+d6k62QKR1Cms/R0jpa4eL
HoBiOKzAlwzD94P+RpoeyrjvywnGBN49OaV4y7t/uQF07xCpr7nGGqWdJ6tSGpA/mPc/lQ3pjz+B
RhFYzL2oymBAQSk03O4w90RvA9ERm8tnBApL2a/BrNBVCmE8PULXVHqpOv45DjdgYPb14HvOlgFM
hiwR8TrWx9OJCKW6cdxJ5YlCJHPzQycME3eKYalvGxKDxiAA5AVQya6IAzlTdgqNojLOyTg9bzMx
R9oAaGNSBNF3E9oocPXbQWEduiDmaZ9v+1Qcpncs1GE5Yp9I9rpEOKtSfYnAkveL9sX2Nh+H47WH
Fx7c2QkLvY8DV8dmvcHFZqq6H5fwfEJt7VvZmseUI0ktMaRx1MPVXButj6AFaQSGgjb3Y2QeH+9X
L2YkPBXNwhaoxAsd1GKGxUipCNOqSe6f868yf72FSqkwf8rnJABJKCsZb+s0dGjljVkdaVL61Dis
Lan8tQhr9mbweEdXyVYVO6ifKc9mcTHSgLg1TWXWyYEyWj88wfjQCs4B3vUsB3ajIFLFXGwLle1m
2Raz7A8z2p854eORaESDKmDC2MUCXUU7wMEziXIc1surhFB1MDTyewCV5zr51I3p7VrVvsmaOWtt
mxcZpvO8+3uttmUEb5O2PQZWndX3VcqkH+JienAG1EioS2N/43ceHrjC1p9lGAJgHXsEdcD1PMH8
BeOTRRDRN9gISLpPEcenPr6KrdIPLIhiB/5sSiJCRLKM4KsnykeS5bAAXRhEFaltOTg9Msae0qsB
fzKS1/VcuUuEH+2k0ZLkzhAlbdZ8IOdBBGL+NJXTiCVYPACqzeVZo2kqE00jngZMh9HeR0SSZdhR
pLch8SBO+fMp0VZk36pNg38Wr5X55zDuxzTPyOsLew2MzuLJs+ycTMK1hXiQnUxDoAxy52erQMuG
QDkIZicm/MKbTcTB1exaysrGsmws3kXnvq/9VjX+yuKiIacSP54/b5nCCuVLf4+52TXlee41QcJz
QImZgLw1FpEPoC3WGNcV7/nfNZsTeGIpe8eMOD8FdFKZ92Yq5tkTRYUGzUVLYyNKUVvMXShKDzi4
+/pACPUBUQCir58ziUzKAXPiTy8KZVwxafuZAyKU4DbFfZy0UJR20V4Y8tCtTS53M05o/j7JYXHo
8wSR6P2fdhmNXgWDrfzZN2mG8murAgR8OtpOteY9r0viXdqhI9FujTJ1jBRBgskPzystT3ZV/GyV
pDx8r31aamSVnZLLMaQYgcnRVhu61z2m5oTeK+5w0v/psRYxntTIzVuDC7RyfcJr+zxxKEn2aebv
y3/KSKXjDOzScrd8ZN33tKya2BMuCEBbCFvRzK/5Ti7dy0eJbVOgjzTALkphj0ohr+H7eKZKHrUR
QjULabUT2fH7E0GF9Rc1oFeaOXnqjKe3HD2M3Umw+o4Hk8p9DMStPE1rRay+xFdJi4oChsmzU6ED
NJfdUpR5h/LaASnGxUZyEo2XaTfDGBrdHBG/1bN2EGwVMUgQrtgab3jeAhfY2tHIIrbwSd5xwvs6
nedNPRK/cbFEhtguE4XHvijivtgoDRmP12gJFpqLUi7LDdFGC/omSjusufDgPeTTnrocVRlFRaMH
cYDAgEYb0V4a7n7mfG1pQErKrf7pAKb2XY5JSFi5+jsdzK30xtTvPKdcDj0hZIkLw3OU6Sgs7KIO
LvFGccvaltwhHfDkVBB/4+FA5dUi9sppIGQeUG0rB2W0e6+V+/cA8dlodcsqg1ieULryV6uCdPj1
ntbyh7nRk+gOaPXC35jwhdR3BjibEZa0umxd3ua3wF5/M7WTpaDUdZIPx6N9CcicIBBsA0lY0ByU
IdV/YDvOB+bg3FAdeQnqvh1y/jd96tldnlym+JbI7Mjl6mm8vhZzJJ6W3rc4QMON6toFaqwE4fqk
8r88i72Mp9OocSZrdXeZnDeqimlQFE2LWSaM4gyJaIx/tk8GU9E8JVz/o5pV4WlyJ9za3z++1p4b
DBwGGAlPxSRDNkwLQUz/MkJaMJgrmSZA42M05nFyBUmCx5BC8bPVBKJPazBZl3e0B+qYy/Z3pCqd
iTNw1SQRWrTHTM2lLvJysqJPGdVYG4WaxGbZjyWyDPsJpsdXcYBU2TIDuUiMZD3J6u4kt1N51gMU
Y5AfFFq7llj6xsBmPCWqOToiatxHpv/iMf30VR+CmXgdtOZycbtbs0qkiZt2VVCOU9kKTsjOVGTz
wvTFyJe62KxROv1rZbBSgWQtuKNYis/IBZVW72BW+QEDEARU2oax3Pn62U6t2J17WUFZ7L+3GxmX
pm3mG78xNyeWmKbaNdZefatIhISQh7ZYLlVawI4sYerWZZqRD/NgQqnW58cQ4h00rhPLKxnd7Wlz
LoqFatP6RRJXsl1Wfq3wKtv/Ue36nvx/G79nUxlzAfgka4p6siLbid8ZkzMoQrfxM0QremHC2e3o
43pDSx2LeDi4mfGvo97JosuTXK+I0tofwOjupH1aYrjROGPkJWx6s3Qv3yrRqfW9hUbrPR+DdsKb
vn0SAMacFn3n/Jc6VzlVw9lnKI9pmLpzsDmgivEaDQLSi4wVLfZzL2CitlVsPnqKgSxJgzlHCF14
Tcq7I8HmVPJSVhCs8+QPcONoYYnyfIISemLAJV7dgYtDKrgns3eeZSJ0BWBRGW2L0mGcQcJ7zVTp
eB+uWfFcRqcgf2jS34rs0mlL+qkB0nbKFMiNM4/CG/KARgi+Xi2g9o5d3pdwv96krDw4qnDZDJ66
05PSY/tyFEiW1kRUAJYSli558i/jgsADx4K4eC1fXu/VpeSAMrkClnOiOuXhnQVnbkv5v55kNQEi
p14yeOa1OQ/773zgjNP5prh/TOKanAGk/1zxVttI3cIjCNuTWyVtsdugfNlOjMJN0SKQaTPymPt/
hJZ1ldOt5K8/wQj8tsLJj0jp+KYhyRMa4+IRuAeWX/YI8vFsOE4piO+O3npf5vk3jkSX0ywnZfHn
ZnHKg0IVOgBYqTDYBQQVOt7G4ai2SZv2NX8lB9ruvTMT6bQQXE353fnUmFdZht495bVE4RnK5Cwx
u97Co4w8tZ1SX7FoSSr72GHthVphDNXe8YS4VfK3wNMWFssAW2Sg3R+ey+MlJZau1a2BMaTrMCPi
iS0+nYXguzyE/LWOKQ+ZX37qFuvq5eppeWRwiYQ7FgwQDfQYDIa9fRi8mzJC18QW/K3rs6z5ZzfV
VRa60rT7StWEb5CuKjGwLrsZOCSFqXEf4wc0DIFCO3jAbtcIl65yUF7VNRnNiDdhMGzGCuV9oRg+
zmn/YSgSZOlzJAsW9F9XlamboTUh3wjaCh1Wwy9OIgRd8VoHndp/mAUFeQgbNV5O9u/EGUQ9fTRq
NRxyJPkpj7cDODEB18V3D63LHCiG5GFECI3+8MhGfHs8XjKzdfQE38SxlIkNqtG+UywGAAKRlC9I
mK/832EqFkWSPzEqmqiHiA4mMeFY2Zgis4GjWIsFh470Z7ZDrNtPzLrfzGASzSh6RQLjl+MBrtMs
HSCh3wJ5dLt2Y+cezCiaCyan3Aypaqau/oemnbglaw4Yjuh/+dNJPeYDVP/k2oIG+fDWv6PCCtsC
0dvc8InaHIOzrZKOfL+3dDiKgrXslHH3xfi8UfZZtoklf3dy05qsn6B7h6F3V1h+QvwcMpG8WYRm
E7ocktK+wCQQ/XfjZE1CGqG0EwZnFitrRMJoGXh/A9q00GbIAbohNVD7Vs8UhVPSC9Hv8jrn87Pi
G2+4bZfgwuDH+LtlhJjk8HeM5GAXAAZrAnd2SZpZqMSyre+wr2piV+Fatz5JYia0QwjCrmlLsztX
+g+tni0l11MUiOOvGmwftByb8DVAR7G12qtVAndftVT0ETBH5cX5bXAr0t0TqwyiG/PD6w1vkXVC
FKa3kRySPkvwReFfUFVuI/qXjTfQeYAZNNL4eGnn9N9iWKRcvcCDqxmag7wnWgivn+MAURSKKlAH
mvoQ/phJQfG34uCfkY6UiFypv4NgUnx5Gc6xAaZHNt3ETReWfe0NryZL+kgp9Adrnr2S0jeE6AbN
XjN7KEiKZsmjfh+rFR6DhBNksaGFdO+DH2NNPPYlbIV6ayuPsmHC9jxzDXtVg7bbdF8kt2qS+GSy
GDLNidAmbf5kGOMGh4GIMpTBjsunbk/PcqnmE4c638v2UdCFgG/dj/JVeb8xgHzDhPjLq3taNRyF
3kk4zLVEYdiLBs1SmobOtWW3rDNTq4nTbbmyVWtST4U6IsAeLb4xJfWRcJ4Q98Q0aIRlX4CHBHsj
Z3q6GUYz1gcygz9Bp2nwjJBRpSYzVaUZQ4cYNdBmhhuZzUOqfN1+ftCe8V6m/gJIfakEP7CDieVm
jlmTNajb/gK4//Cz+B+00yo+AtGd/BW68MnpCA3bbiqKR9mpKwi+zwJX8WQfpw7DVBcTQ5H2V+1H
keVmsdoz5Y06X68788NvS+54qQS4x3KbyZ0cBFHRBYVXZv6QeS0ihamX15WMVkaFd8vlhZBd9mzr
oWw2uLAb+sI48FUsCOeuHTYfxFShlYiiDQ4ngiXuYXvHq0gxz20NULr1uQCUocCbHuCZxE0o5CMu
rO6kYWkXqFgD9xiPFOPwkz1E2FZwjFSlIm7q3n7bOMuzoQoT7GCbH3F3xQ3J4wCxcWStKwA70zZ5
A+1UOuEFO8IKtR+ndxPVzPxl6Um59ZNkt5hxu3jaIlBrf/5PXvDE9FMt5moDZalYqJPBpgr/Bsgk
dPSHj49g4BmWgTB3VqluJrhP0Mbh4ii39WbS0fBGWd6ZtjxqcKB/Sb893xNKg8jqvNVAPVN5vrCO
wQ7alONRy9su6i8izWcoN2LugnK56eV1JosGFti0ZJfgCIOy2CKMH5MDHzusOSZoxThQLDf81M0c
yGlMf3OOV1sRwGoZdjDkIL480ricl1DPnT42SueaEjvdSZfQRl0J0juZsK5N+vKFPHol5eAD0EB1
WCXr/ZghYVuRhRpl2caWobDVsGun3dxIhVfGxu9fjv0278S2qwSBVlS0YQZ6tIQllfNN43vD7qVo
pMAP7mVd7sD2cuiyu/fobD3PCTSKBidLWAhU/aEhNgHjOofiJ+ZZoPmrHicFCzcRVQb1dO/xwuxK
0F7qh0lb6O+m+VwT1kTXCfARo8w2H09D3kEbBl8dJE7Ks7aPfPG+va8ByQ0rEF/403I0ikd7XO6w
uXEhQutXzm3rWi+O/sW0jblzCYix/2hFo95TTuG5oc2zbDJrGmCp89YMBG/otyzkTSW//aA3mp+Q
ClNI6CVl7eb/Ku7ZcJv8/SHQUcU6b70As6bkHe+IqDHyq35hFtLwoEUPokhHFpFylXbwrVrYVsyz
zUrWKp6cCiCjjXvP68GJAMIzT7GiOysh9ZYIennKp0z7xkk4C8vR5xp6QsQwcYPtq26Sh6fwS4fX
+NKJUN1VNAIJCsqmNV0XT4UNrCxUtLzhG3hvhbqK4RrSrKHIbmOi0sdHx6rqwTZplW5CIiGXMF49
GuZ3zxLIUffKLK6MQLpfxPkoT3ne6yoNKD52a2NyDuuQU2snbKAUmkPBaVFAd7/MIUYpatxw9sQX
TO7DnLtrE73kiDsJ+3FZC9SzjJDEQr+Q3KTYIqlCBj8kfkDzhdXcJXscBRRcllyDoH9rsI2kCoBg
VcajcB+R9sJbX6X8eDitfyNIl7/E9nGPBbwwozjoFB74J3cTOyD4+9PPYbrwKDtzmTJgHNllHXoV
pmnPp9T5VL++AT2xgcCy/bPFB9vic2KOvx6/2Zy5jy9ZNAKgAieKVx6oTRN5VixLE6TMj7xddt0I
me9fb00Rg9sixYMayDW0uviAqKP5kEbPKHFN6cLcra3MHm98O6aEhzuDA9CKcPZcPbxI4BkIBmvU
A32jz+FkfUJLC7lIjSMToRinC+QTkuU+H6zs1+6nWtiJ1vFiX0UAOHRpU2s8zCj7mAobTo9oHaYW
FL+Ihpp056cAtrMxP6fRGDcO4H4+Kj3CkNyQEc5n0GVADgXX/jZcaOGQv3qB7pakv3RLNPtyol3o
89023cLPT+FLuOB4/RnzVonyaiBpyLupsFOr3ZqZb7vcGQymQ6myXk8hDKgzh/FoQPnD5SNwDZbF
WSzqELg/QABL1EVj286uk8w16ZeDhKr7yfbe29XKEOBtDQlaY1sGwMXaX0OOHfwiZa9Lfelipb94
6WnUaAVTYB0IWlmbTvjyV+2NCDWN8kkdnz2KQKsOsu6nMO1k3PKzy8bMAaRMQ7lJXcftHNl11mK/
EcVhhAJd2NGAbEOpflYuT/VZE26i/GQnfH1FBOD7fCXI04RZFwONBrCoug0aNH9Wfyob11baiOnQ
rz8srpoIhJ3QG7boXiIvCg3NVXKmmu+Z98rxG+CWExRBmC/OyQMHXeU5VaqjzsBAeLUdi6pOam/Y
njTaH2llPieEB+MDG44sNGRNzo5rvNsWjP7yNF/K5Eg6rneSE6mAKMlt6ksEXRsqKiEt76XZoTDc
DJmZ/+G92kp9svYHMnl2XpgR9fkxQgRBhTjBAl6H5gx4OQ78Us1R0+uVjfu8RwGaK3awwjjjrVoi
cWB5sk9BflWEN2abEh04YTseYrgLAL+CpQ7coJoAxJNp2gVmZ8zmp2Qvw3bMMzi3iT3wlWtJ2bWQ
8vVeM1wp06IcVRh9MvnRwv7URUhyeCH6f0AO1l71L1+cmaYpSx9s6RvwXxr2UVevHL3Islv7djai
i1g31R9FiQf1PfKEuu4I1h90biVHRGMrtinI0sJFOBAicv0pQ1FwyqLqGNIgWNBy8KGzsHXKiVCK
3+B+PbMu1VvJG1G9tNfjvexN18X0pixuAgYsCkXfq0oGPVGCWIWz6gjpcMm87dPBJopLy2eFAnIY
rHQeuScG10w+46c02zTnFgbG6NsSGjN6sTDeB5XyRRddf1NzTJkHsunlY0Cfq+UgL/ce5ktHKvL5
saboO8zdGm9nDHLNcQKhFARYkWL1lz0IkCFBwGdvxxQAJEVrIJdfO1I1dtrKRG0RuD4Tp3XEztyk
r81kaaJGKRC9R49JIKnFkw8VCxJMsGKqS1mU8zOdxy5sVvyJ/WSgwaBTeld7yEu7wSbG/8jNC1ej
M9PkJ6p3WnrZgqXlK5AKayfyIc3Z2aPlU2dY+ICbiW0TgAa6Uc4I9isHLBLbtGM8waygk13CRTdh
2PC5+2KhE6RfvWo1Pk2SN+/xAb53kLsrta7LuTRIrUAmdaz9YtYFks7XQkIjpl5KpWMcMndD/MHe
NM6WNv2/UtLLdPVbzR6GCDFHjiBM05QzjXCoHR6gZY8ZTsAM9PAURyZYBr+IOAqE1vTLg3d3rEUc
T630hgxBuQzQxtgdGCChvljZN8MHfI+jbClvT46Gyrx3jZHi3AzRJv+f733NQtPRXCw9S/ilLPm0
3WgXwuLBzQwRcsqb2rmHnaSeVhXeJKBMHT+JVZFk/JQ1Tr0QOFYL/jpdAEnG4hG7dLvXnaVKbOEi
3mimWTYmtMl8mHhL2Q5Jhc36niZVRyAGN7Kd7crkbVeP2uGj50aHzb70Yj8OTyGWeAEMobIkERMI
qGfPd9ZbF5GIB3QmMFboUtGcra/RhHK2NNkFeuwC6jtcjyhWMgxbsGt7Vt3vYPtef+dBHZVvKOos
LwpJUI7sNFZviZ2OjrmcdrKVV4uBbgPGkYHW5+1Pq0HEkNtUUCPN3eMTlEr4h5OlZj0COkumO7KZ
f6Fea9WlxTuRIXO4qfnodfhRSC95sX6mPKLeKBbK8tVcHqnUXExPiSIfHVjexthbTlRkCdWj4DUr
CxVt2RQUF8wgF36BsWK/qIPQ7aZnzrdvrgfkb69vYDqdZLYvu3dfcTb29JvJ79MTm0OBsE3LCr66
zBjhdfZ0L9B1oiQLUivvy1jws3ZuIK+gxZtzVN6uAoBxZQVz4j0X6lBeCqql7LpDpNLm3SE8VVFI
vcBE7Oov2gw5fXjdH8xXUkb0b5UgHo9853pjM+ovldEk+n7wino1NupDxInT6aWUuZPz2zbusA1R
zpyXNUL7kUJ5aZMh8WuNJsYdQN3Mnx4kfkYE/8JALzV/3MvVR+5shfrYjK6rDqjQF19GcepKxG30
P32oL8Zdf43OluakS6DYp+r2C5+i78pYKj6ML5FfdCGsaYIjvTOv8gqxDGMDHgEt5QP4WJfLHctt
jXfSIQZZWS4eDI2i/NMRfmORFOtDQ+lkT+qu1JWf8aYzYtwgfD3UKinW6bVoFAZCPtN2rRMVhKNK
7h9iS88IDeAUYK8PkSi5OJx28Wth8KipQB/LZhB7XFcYCXGCcGCOgRAtmzPvEVvaXB64eS1HdQ5l
37CE2C1TASlhUlyrVjxJwyqj7dkyM+blxnc+gQeEEznNL5zoXFflysNK5xyYw41aSUCV7pmB8k03
ZgGGkaj/XwJxfHeWxffLNNNbRZIlLaOuo6vgwC7TEJGmctNietC9+lGNI6sJdKF0W36b03BqMnUa
CeFHNKKfiw+gYvsZaCS/YU2cP7LEdK/9NmBdcUC8D29RJqm3Zvqi0RlwPM2dZyRC8dI3kanycUPb
Sxin4tpaNwnC7UMSVLJpsxzXvFfYZTrspuiEj0H4LiZhKBBNYaIlR2WUOz5XLY+COLd8vUyskbgE
hpM/yuK96u3Aq7FUaEqsk7va8pZU8Meo9veYJ16jpUAndlMslaE+LOpPCCTpFSYa0jIUPPfgb7ND
J8gg2F9Ekj0OgmZvK8tE1AneBjmlhEy1vLODB9b0yThRl5QJI1U5hU4o3VL/Wv4hDl372ZuBs/da
NTexWrfgu/OjRg5zfCPP2SGY5LBSscXB3BK/+D6puC+SNBkL9p48ORclUfPM6ZC+8uUQ8khevBn2
KN0ASo2XeuLjWVsPEkTwAYH6V5+Hyjm0wWRpUMZ9/FpOMnoV1CVYFOZDQCwu5Bc4QyU0QZkiFq3I
BVaAl48MbkjvYKgXscHvldCIRVVT2ra8lRwZO1l36DG5MUEllQqB2IbEUO97Xe2VVPgHSEXWkPic
dUpxh6GxHggTA9Bvrqy1uNc3hWhhuTVGU2R/pGVGQM7zUL78Q73odzeAsM2YeUo7KYfFbB51SV+v
XyVXBMGDPnjs85PyXc8uBAc0Mv3tkiMrZAtnH7cU3ouD0MBje5gSUS8CMgtnkFeHiD3F6D6aLLXO
0QrZcf/0ENC2fCASZCSo9p6Tx33SInFmvTVy5xxe0CJSrPLe4holLaStQ1ORWjpDnHPA+Aw2FPCU
n2SLdausIzweE+ap28ffu9Qj55APi8wEb3Lyj6B/rNf0HCATveZakCYDkXsb7Nfx16qSV2MqeOXa
nN8rUOMLRN4D14yIa85ZKsz/MC2Lvfa57ETAzYHig3nuhDOvphwprx2ha2cUiqQ6cGgixSz2+Qnp
IcWriFrAmYUY8Sd2MX+++U5vr15kmcJ8fvtms2cXefxQW4gn6aG8buy4ddRt/oyyJ88RKDkP7dcI
OO4MZPWzTgeT7orP/Mt8jRx2wvsvPtCOpCG9seCzOiJjx2O8FsICmln00NtLwSUmIR3RNnuIMOWQ
1P2joqbY/1Amnu8mABbtzdehCK3Hux8oZA8HKeCF/3xwZbz7qylZ7LQKuKS2/MM0/j6qyiJvvbn7
6GFPsKPoXZVHdzx/YOD85diDGsPVALrBtoop0sScXYYbN0bBUWcGleSEkJph//VQuVd20hYF3pKF
sA0VDU3LZKm9fQLRugte6B6OlSwJE7E6bQFHBdXZBK1IJkCH7z32DiKZGXIBN9LhZNhVNB21Sf6l
tzW/D7Q49SYamv1UZ7yDKdxrDnOAuY//2syr+0ly1KVQOudy+QTiXJl8TMi1FTDexpUzbvXWN0EM
GqzutGxD5hK5KWT1aoFjnjKwSizcRANJW/g3UBTTkBBQoJSAvTJbbDAeZbjdk4G37Fvo0eXrYGMj
/84cpHLBMtkyTkmTxTHtkMO3XWFw0h/71UAVUCogLJyVRU/MstNYtMIB3Pie8wRVbYRuTU987vcT
J8JvGe5t+hO8eS/evYbDZCorY/1JDkJ5eCv5gmmpulZpgwpo2Zl+g8w22cjuthlcWDPcaEBfMFhi
2o3P79wyDEizKUsZ8Wy1Vh8wngQyLbP0ThZjw1Fc4jwUGEU/wkXRMLYW+UwYHjRmBYxi1gUeELmt
0tREE/NvYmwKd1fF3QVdtqKPqtR+8U8YKbWyfLioSltVXuTbBW9AjTWLD5ZOncCv6szUfe5XJjlf
ji6JiUeV6TpLeSeRIz57OiChm/ET1PMS/K4J+CB+I1Oecy78Xn1vWduvTW6+ASfiYsusHs878221
utSCngecPqk77xU5vv/m9fMrwlyWljplU2oj0r2VRoXHUjn1GXR+GjZde8M55YkFpxh81x3K+Yde
zU6h44TWbxMYyYyux2cYM9og8NadqVFKAsWXlsOIlZlGJTARZimSkZDuEAGZ8bGKI84DRKLQwPBq
4+s5GlLXm9k1qQGxv6uWBI4jeXtu/NgX8/JdLreWy6TkmOq5LkV54OqgS51r+yN8d4qvp3WVwp39
qYGGGVR1d3d4O2QPuRK+sXn6Vd4DgkipVuSO/vGyvLuwp7sZLUHYbnb3FP4xYKovGG+5U+CjbPxb
3BqJIWI4oBaOvwPPyPFnweNTEdK6ctKgBybOJRvBPPvAdyAmY9owCjMADjB47UUVJk8QLwg9iuDr
LhJ8ccRVnDfIXUaoJNvjxamXQob95OsPoqRFzqyX+53y4DTL2h2d6fNtbt0xmDrtk2GGRum/lwI6
ASzHOkA/tRxdjEC461bWRmyyxciABfTWWh8bU3ZCurK9Or1f5AutF/H0uiDfXOtRTTUi1PVEqcZP
4rVy75cK+GZ5/EXg77D9M84Iz+Otu8qDCM4+Y50tVhLwpIvH7+mGfwpBraemntb7frcEkmOEZHki
HEPD+o7cGe1qdjjeW4J7Abkwzg3hZlZ/l77y6UZuZVNVOCmBXP0Pdfp7ILrQKHokda5WldHuDzZj
r499zthxFnTyePO9RJuPcxazUZhpAZHi1EcqoAX8C4HlLOJDCdQVbAna10Lh5S4Ya/gTfo3fovLV
GHGYVcMXQFl4rdLxtMatgbMr1daXLq1GioDmwy9mWojGZQXCVdu1+0mymF/WngdbMcZen1GZGTJ6
zOoCfhCJcKpvD5DJ8ShOS8thK8w8u5RdF/vUJ5ZMLEREBHImIBL/vH2c+vlID5T5P+Z6i8rk1/AO
MNYITgqqju3Q+0Ws8nfZtdzbOln+Dy5Zet11E762gnrxKWdcqqRrQkiKO548xojk3SZkKWTnZHX4
WcChZOdXW/CpSibWbM9XfNbLK51jlH+hlC+pmyZ+zlWitB0sFWMyoEz2iRCN2Sw/LSnriBcbleQq
E0IVFYoewShbDzmUhP/bXfbjMUWTdXdD71mcloXluLCSBeGnrPNp+GdExW7B3mptBIVLszr5hRCR
kEAn2tPBUdV2WJqhSPh/zp5MzZ898i6dN9NMWaY0YfF3kBISuIjdnOP5l6xA0XAcyriwcj4+xXF3
/0o4s8EIc9mSBftzrkXDJ5RzcYKL5mGwP7onSLoJXsJ2imMUBquWqDxr/Es4xwmaEwaCK7lT+1eq
W9r1XGvXK+bmbKHjNK3+pp/jXvozVDNM7hrKSkSTIZGBGF9sKqPlo9wMCPF49+6cqXnZ+mewTnYv
YqxtfySHlmmPsEkx6lks/076AjgclwoWX8bVGOUZY8wlR784oRWzUU9Mzu3g3YhplOUOJCT8tUQR
zmKF4nbvP3z3zodKlF0x5iND6LvwFsKIZDpkvj8kuYmqwi63loByhS/Pjjd0R7NLtlkFSUwQgOgL
y0Cu50ndYGiGVa08JibWIZoLNw1Q7p1Ln7UA9/LTtFvSN/hMv06pLzBoRuiseSbDXjXDiB/zZfqR
iQtUiGLrlFOd0pqQ88sJchHmBDMR+UFkFEn1X6c+M+mf0OWGeMkLIq+OGNFt7Uk8vpCGh/477862
l8VmFs2hdzdONeHX84cHAxUgAsvIg3OZaNdtwhbGzLjfEHaNSIU2ZpTtFPVG4E7rX+aEReEoTmUE
/3gAnz2tcRjwUwS1d2O0SX3Poaf0G+EhjyR4y+0Mdm37nY6gIesmQRSX8GQ6dLCjLSaziTgWSr+o
wpns+Ue5DrqCJynhTOkwlI9d/ahj45qZ0omMrkkQV4GmhTagtWVqgXkbPv4cXN1mk/hEpS/fimFX
+F4hEWEHxuG/84mw/vm9rKOfJS7qUUf22JcdGK4V835GiuMU3QwJ3mCvXel/QCZ9GLKnyYPS711O
4GFdQcym7WMICVnBcSQWLVFGouCryA34wuDCm+eyBYN6h2C1EtIRYHh+ivZro2shVpArdxDRVssX
xHEOab1bgrEmT8tzEK6C42nl2ms2ELmzT7aiUpwSAbUeFPt04KkbJmR5C7q4rkq7b7LMD2grc6AH
9uWHZZq0mGz2pLHf5DuLFndil+twofqPAV+bpx51fekwq9DP0g/Zb1ppOeQYHKBIwcH3GUE2ga2n
AssF4GIQr3yf53uW3C+5y5WHm0sVNancyOd22zwd80tlnBhCmGgmjtzDHDADFdS9o6wAEdCRG7cv
Tw7uQX+JGB7+VbfKHfnJ0EQ/lNVYuToznzPKFG6I/EXrzNLmKlJJR7wOOj+R+198s7TVK0oAAltV
58uklOdu4vlhRXpkZesxQCVAHsLdYKt+9kJh7k9jER68kl+5iVhVHW651we/XU+PMIEhBoSGz0c/
Wln5Smb+GVx4W18a9ZNNONEe2cbrWJ/65Yi0VjCU5YHjxki5mmi9JZtU0LGfRaR5p6Q7avjVJAY9
evafJyNPfUsOYZpv/JrGRTC6XQJqEwSW6mXMG6W10uUMxv7Wq3f/hSP3dItLY9ROxoH7K3FwMhve
uf5WbGgB7TTtir6r85uxFiIw8EvvGUySGY5Y0I+tHokaPVqUcWFheHcJEu62sl6xTSrR3FpnfKY9
KJW0sRw8qUHK6BG/LM07nlEdS+j1lUJBFv8qg0DpLKbMaziM9V84D5ctqA2uqiaognFfJ+ySWKC0
pfIKjBf8FEEL59i6sJV+HIA/k9Wnts+XBuWW/CILf4DgXXq371Zl8y4XcGvzDMQU8qDcbyxRbAMH
c0zJv53XxkodcdXpyuVMTalvYs6X9suEC8iSYcVxV0JnOBhRVxlO6e56hPK1nRMw9L8zhq/8JSDs
Z278Rm1IXAYTZQY1yRokGr1/8dXh715jznfQBlnfKHTMbD/PLwsHRzGBH5iq/1y0QVYyR3mdmamC
zQ49XxmmGOg+i/aj3ZUm2XrICJsY89O1teeqYjQjjHIaxCTNJXiBHN/sTlc1J7xT/YPHiSDwV155
2pVg3jSzy6/XNoU9nkF2gR66M1Vbb3dbHwjr0MsLR398YuJhzrmNYLE9o5v9unAQ9oghXCmjpEUT
W+pZhgmGNhjRFl86ms3WY1PRfMkcRDmhZJ4igCrN1Eb6OAtpJ833dpuA/1UAOeIDRZNemjNRAOu5
dyq66CPOcCC+ewACknwICYHnAi3mQJzpCaFr+mVaQnS5kEBo4IGsc7WKrlJHrsy3yUnqTqaAlbYa
rYUK4kq645h4CJvmrZgZHaBBHrVYI1hf8pSjbovSa8tABx9imUG3MaMW4WkPcm1wkIU9kyCWVbBb
NYyD/Xe3c7kaniJ2b+DPSPxhwf1d3JV2/a/qYhBdXYuOjyphmCRZ9fe+hBht81SdOrmOzT1BZgzE
FM2l7bcriKqNi+VwP5wxsyMXJBZ272tuW63Dp0Jh+b0/AR5q9TCSZVyRtV0mzDCOPWm9Z0oJB2KF
Mr6BrmtARtct3SgSjZpe9SuDS3i0gfiVI6n09QbOnxIe2t1YMA6XGS3GWkfygnNZ3ZEFegkfXzEA
8WxCqyyCfS0eC7tDK8JH1VTw/nTSKGsqu/XWw/l756JQk+R3HsM3cVuFgs0HTeN1IJRdeE+7Gii3
45ji/aWkJ41duME2Uz1du5wvxuS5YfV2ly7dNjbc6MYPy7TFfCGhiOpD2+y3UOUZeYgXilxaxjPm
RMocwuuBs9zg1vtGXcr6tIMDWzsugoJ/K0kXviXrB7bp4PYzVJKeYXQbC/01e0h51ipurB/FUdg2
lmbHd9kbFoQxkMmn/+10cLDNjkhz8y6us2drTKUqBI6bWkmbrCEwl/G9jyOh+sOAJN4oD010Crys
92LOQ5h1Fwxk6KBFG8rLlI84BV9Sb5LHieR4u+Gfjt3HSVT2096DKiMxBCELjMZjOZYS6rksZfLi
M3hBSC/2HxFjjIGNdI7j+zWv+XQbHarYuAd4lgiGYME4BzEq+bS8uIHusbqkhlCkdvBKeehvEXpt
9DKnkwUjduridMTz0bDDSp+jBdjG3hugrN/eitL+vlriY7UMUQBk0DyTjMCTk4aPqqnSqyElo/uh
VJwXtASX4eppyXZSoN3/h5YnUnZbgyvCldNliOuRvHMG+Qc0Abg0pqVOmpgGWli8K/rtu7tOLXSx
xyZiEv/LQFXRcKpxG0OVxft36n8wfAr8F6P4uSkVfQow2chdOzTg1wGL3yiVnECth9z8PutDNwGm
jCLz0wyvsIeeBwxboq0H4jHldkCC6l0b3wOzifKtdyBZ3YNd353UhQqQ3J7Rm6+FSTD30TbZrEs2
/+TJX7U0CbbbT9Rfh3FFjGiUlAkeBTSx2SbAaq3Fu77xqZO3kfzGA7zlo7SQtn2+1Q/9+xNw737o
ndiJ1Trtu+jJOWKGOFhhAtYsbfbyMXoYtV0+rVjvCCOwYKB4TATVHwPvFBSKYsyaeIncJ/H2z5x4
QumfH5uA96bZTix7usdX7qKmexjb9lBtZFXvw5CRMsLReF/xepKEZ9q6DLHO/srA0jPwvhZZC9fY
sq5XnXBhqdVziZJth6I+hMcwD719ZXcqvs0yEbPoo/PV3xy3ycBDuld4uq5HM8/D+mBhuNvqFIgi
aq3+pJFkPzHkhtR0RMFpd72UE0/vtjsionYFVpmYpy1/Nk803IOWOffdEZi2XWw0ZoAwwdUuIgJ9
NtE8YAYVPYXabPRFp2yBIay/2i5TX3jeZjh3MAWyUEir75KQx6iEc2ry6fwHjBYRqbDsG8sIomw3
1U2BajSuts4yTxbEnzB1OUxA8QdeMcx9E/FvEBy4Gz9MTpJPjDowVwsWUiVQbRf73M6dIriVJOUW
O8dSmaBJOMCbZ8pWP49EEIZquepKEapi71OiBxcOompN2beNrWxlGkLRaOOgwKu3Jsc0x/7xtpmz
YvyylIlu0JzV87NskETzQozL9hx/SIIpUg0pYcMX6TeWCgWmPNSzEcvT/uMpVtaDuPXiTgN7/ZKZ
iqGfj08eK2LmwdiEgbVp5gduyWL9OqniwEW4w3LfthIASVyevWauUpwoaVRQTYcs8c0nq1DZcBNe
7o3UjDwQpaZl/jrwX/1WcLWjxOWj4PUdss6geSnf9WF4igI71AtF/46M1j6NeBulzSsPZgbkpISM
M/u8P4vzKUylOVt3RV2b5w57bZBwpQVRVD05W8J2sxVgGV2gUPpyv25Z9JuIqZCLYLWEJEkhnNQW
3jdt0pEghy85toSxOkLypfTGag2qOhzZDTW4akg1z3/vIjpj4/+H1gHEd0LVJujwkuRtY6gk8xcP
zltFXn4FPeKFd5Kavl5+O9iFE6ONP1vZCPneVZbM+snLjrL2cYqediiegKVnmYF+7XVgUzowk/bI
YHYRldNYRYDFT73o0aPYJDCg+/bvoM99FvtlUQnElE92qgSntm5/a+UEE99R/YWGOwLY0HIm41gh
BUrIimVFTZ6XS1Oo6rBFP87uaqEH4+0pxbOqAtQu9zqUh4OiJHaVZzpvCtcCNB93MP9yf3PgC3iv
lG6acS/LjlRfLsuNubdbdVo9a84cGO2clac8rh0oJd/r/J/lJhndsQ+aaW6qhvW34gJCe1tKVGKI
wc+vrZ1sPpk6kt+gds2SwKTSQjNejyMbjXHhVuQKn/LmTywIDpn90yFJaR1DOfLdKW4DbupEuGTD
sxL63nUTTD+by4SUCqintfDd3JLXAybmyt1zxXJVnMmL/VkRRs4IpDaO3UILrPOro2Q5Wha3zaB7
sS0C4qkMvfqpgsirR3a/NQoNFeCYRUTSvEdr+12MX+L/HyVSwzbJIvuUqKNJe/XATbTGT3hb96uV
/G3mEHW/jgjb3mdlgwMl6snVj3yjiNJyMbrXv00f/3/2DmgYNzfY4OvRLR6RsEnJGG6PHZpFFj0E
tV/mtYeBFg/TxySIe6YpdmLjgMZDMQZu/No6gYf/wYpa3gwQspwzx+0pXULBT8RB8CwvhFDCy6Rn
H59pOPTPyluQ9i93rmgzytHQ7mcTOCAmiKPLq+kDaUXlJHSYisjZBHmMKh0wILDPXNvvxR9qMqhX
llDOUslosmZSemlUNla5cg6xC4vVzMkXulKdKoatFbne8z/vplynpe2ERAd8Vjct/zU6IoOwmysg
zPvnVmJP+fF4+k8ozhctubcbLO+Uhaw3CzdUkF9UARkm39zmnFf/TWRtY/wlxufSFY2gRUkB88MR
Pt53r3S2i3mbivxe/4c+PjR7MluvhX5enpCtqxm3qNZ4Tl273eqM3dR4qFjffEAiMcB0b9Kayjm2
PDKvXkDuKq/uYfXcfJ2o0Ru+fGPPZmEB8jWDDLZO6YTr6k/4Sy334FG2zQPSC7CLkV6uOKP46Q3L
htAhu4RcU2LT2qBmUi+Xp9SUIR4vR0rMGo6cLWVLR2wfjB19tdRZ3XzS7aDJ3KuWC0cSKt+5XWoH
n42ePE0NmbXiHunCHzEUpkauAzRSynNYTfUAD/EhS9mXnM8wRphXPVo86IkVbo9LvxgIJnZUEuhO
OmMprD4PNsqX6Cm+xcHXZKCGGaIFjV7SUdns7II4TAhyU40uBU1ceAMNTLXS1zQ0KyO+WrrbA+Hk
ff3Qz+83iL6+Xl9e2xR22pfkwaUoEzprl6sKURAv+5v6VMJ3t2Cvv9k42FpwDLn5w4rmHd8gw+OZ
bQzultwn3VqHTy+WYa45vw5uOrQIaz2TB1c9twa9k3AgSsqymAa+5loLxGl3/fdrZL4oVG/c4CP3
B3wkhrm38q2tgz9IaSQrsoTJXh+8houFSjShEmoSljMCWnvolFvKaB5zd09ID1rN1SjEPuKOqJUR
eIB6cB9emUmTctNd7Ch0Uct1mHtH32PrZOHG2iLPJNjFOSxmLheQ1m0QZvfcB5aVukKMXC0/s2u5
NzKvCRpr59ieLJcBPrbOa5fR2skOJK6D5FBfEqkrvyHFdFwQ+T4QKSzZas1EE9jREDmkhg4lCtO8
1zdS/nlAP++uctLEaidNK2xhGK107nXshJCzz3IkheewfbGZvo/vN+68es411a/rIaTzlV+izVx6
u3HSkphEVuP2OQdWoIcqX8TPWiBbDCHSvcjmai8CyJJv2ll4dEkAscc2GBLtZf+Gf/+osTiowhWt
DVaY1S9GnxwJJvgis4PVtIo+FXpq+NqlT438lKXi1GaqiNJ5A5uGaawweiadwx+nYmokuHgFR46p
YLl/yD+wXeCZQjz3uYjd/aa3UybVxowkfu7ufJFQeymgxP7bRrbuyKSRIY7SOgxTAwX8p9zXrX61
DqT2xw1xMb9LKl9XBdHPGMN33BZ6nG8L31AcphL+a2n6hxe//aO/pFujDjT47qmEDT4EI/gridMW
GiCYgiHXJXs3z8vu5NPI6wvC1cM4yBXklH2CD7evQgD386uspy0lhpX9LjJ0Vvi/i7VL7JSfy/BF
4KWn03USwFocI0H+ufhVymBA90AuDKF7ewT+lilacGOodG7ry35Y7D9olKiJQnNbfZ1Ba058rwMm
/8lXO//OyJdpnImMhV9DpmdRPlJEv4lAPeaUvMb5vEEbkzdIXWmPpTpfLzdtPSZDdt9yCYLjBzDq
cHaUAltY4/3JF7Kp7CQgtYMqh5tqdf6eUsIQCwPa/44h2vJPAXGeZ5NKDYfmStNBPpmF4xOzCppz
GGVCi28+PcR0DuRdAswWirVvJgGLc8l0o1kW3Q75846SD0yhh6bBO7QeYHEHFOOMe39p5y0cIWGk
gjR0b/YD+ZAd97iumPrlfmdBrJiIPmZFVg21VMOYBtPiQ8iq7kda0a8vhTGi/ENj4E565m6z2rca
h8ND0dvfwWmC8NAtdkmuCOZLJOu+6xetDDf7aU7Ru7Cbv2H0tleBGMODwId/VFjkXuGpnPZxVdRp
9h53wX7BzVTS094gKRIfkoELt6+EFNsGkN066eBj2dRXdGYkpuyL0tJzzr38iaMjSECKktbqTgRs
a6ltJNvmQFCM1pAtOpJ4jJeFAFqfUQj1u38mllsF9MaZw5SCUTTfcvqeruA6fMkPd1690w5GjyKR
9P7i36m2QCdj9A4qzAJ8zDtLwM+ipRv8OJCzJBantr+/tqNWY+J9DXWTIS2VK3LwKg9qtrVDjlzz
MnfBzddnRm1UZ7Yb1808YU9EZJNpuWBvfSb/Ha/OqSX9SAWIErV7tTqqpnBdmbIg266zupaFdUJ7
xr50PY5xx7cA8RFKWDZOpv1tL1dYEDqGDQ6iXqmlzzj9vxQcorAmfaPMVukBE851VE/UBFp4DITf
9LxrjL9qAW7y31NxByw4kTY1MS8KwJ1tQpylE/OrwGBF7wgTAcGiq2iss3Gl1NrNsXS0dueBDxpV
rE2bYHec7Fa+1scSQtn1wlrEt3zBpjnhaFlpSZ+0wAl71cOhqnoO9F9jEz/Nt599HX9efRp0wius
304MB970ATObGCOkNWC+5Zjceq84c/HqNdf1TauQL2sHM08N0V6TREYAfMu1mv21MZ2EQf4M6EJl
Y+vHsm+wNlb9WDu5sRDGvAF3H8ODO3p1OicSsDig2uV0JgTlUeR8gtp63xPdgF8T81IkA+gUaXUZ
ltLtiXMbJ0oet+cdLws3II+8qmN3Mof/YfTgbAYIM+uAq0uZcaOWp+nE55JgIACoQgelCd2Vdo4Z
dw59CAxFF6UHsZEtc4dzBdBGYUm/9Uo9P2x3kavo2Q52jLm1ilg0cjniTrwkcbDEdR85tY7+vT5H
Z0S61ymbk43LTD2hoyXWzels6rf6FnAZigHznQphIgMDvI2uAPhkkSjwI4XPCp2JxKTHgWGPZgwl
3/5SjuU7puNvv54CpahsBrPfJrEGH7cIj7Meu2eVdOIrti5id9t7S+5eVK7eX4MtRn7hjYrwpyrU
Ftzj2Xrx4XXwf25HwZ3V1jiXsASgjRWsFWHGofTfXQCdGr1nGtQDB/JrBzYwbHROtCmHFtb1PVFp
Iwkl9gAlK7A0mBA8hcH/aRc9jBTCE0jbOdH4wxGYO3XZ5m5rooyNo0+ZhELgLRpa32v3jbfkLyLL
xRbcPl5BDCOr5nHr5TB2zJCa/Wfc8WnsGCWuZh5Fp9IxKOBQfHC6F3Oxt/vAa3FoFIgfHJH+m09M
xzjQ/221pzXV8GgKQ+m1FbUaXdEh9wcFTwUvfq7HeMdKIdDuQL5vcOzYuQBu8uVkUKT+Mf7d5bMj
boX1klL+gPPnRI08DGuQQV2pKSnhQCOC+aWIdn+3Nm1O+TBEvHaPZPf1tKbLS/GLGFKNzZ5r0Mfq
nMiJLOXwExheNqqph0WROJ713MS4NSMu2WpD8hhjO0p/82337ABXdb2SNFRHuTdQ/g+LEsZ8EHuE
8kPGqpnJsgrTIfQpNV1ybPf6YDVCEPAzppWSrFPUfs6C0aK5hJx4VEIHR5zIhKNLBiuPHBVCN/bu
exFwpnWHClkmi6rn6drBGRvkjX6kjFuT02EkLMtijHWqnp7Pr26johvchyki6uQhqs94MxJsXG59
P5PA4Sc+MbhPg0C3iDir1SFxFVwyrd4mBEbfoDe9em9DTs5e7EMDZ95IDD33md7saBhcMpbcyFgQ
x/CCdemmsbs9qp9FaGQYxl+fo6L71YuR9R6eLbmSWoG2nxES9NG1TngRPRuiv2sz3TEnSIEtZOJQ
9Y/mCehM1SJ4hZ0QsjP5eoD5ZHao+I5RG7qMCzW1sWplvozWT16Q0u0yROORW9CRNQmfqoCdWHHf
EWpRyLrKcpAlodgrizXwVe3nUUMs1ZZBDJncw58he2p92gyPC86mBHU4Q214Ra4PwqFeDxvdSb/j
FKBWPeKVJ9dsR0WHnOc+cS5Ymtnw6jEMcR9mxo8QLCuyZfkij4KcZ+RkHhCDb0bOsLb47cyUpi3+
wu2pMmooqEwhAs+7kywaFw5mMdrWXq8QHEBuOMoVGQ+uya2ZidrrFaOVpHnJYLTUKnTee9ZeOY8I
MePQaqdcm81DdvljWASCNJtPDQEIrsXHLR5ucBWXOyaukI4kv8pOw3gj5j1XQaUYSzsxWCrZ+1n0
vWcmKwzwTflO8uIvP2cWs7B8a1u94hlzWd04SAY52Qv3vJY4MEH0w+1LbTa+ccnH1lYAQJpZzoWu
VK0FlzLEwWal+AOP+KR518V974Uhjp2y/CBRdP9YI47VVtZXuvvSwbWzeYnlii6sUOrPnryUFk3E
GevcrS8CHbkrbxl7wRa1VvPKiHz9KZ5YhcKX0ZpIoc8OjvKZAj6W44N80edcg4mhM+SNLrIliC+T
86O2alAR8JnFdl+cNV0F8CCWWgfPXomXiAXSIUgCVvf8EYCJFr1lkM9K/hB9PDC4Pitt69hDGuMh
86ixAXbf+mYhA2I4Q+eCRXMAzcvS8qoawPrwBJUjKsR6sW0DRrUmQ6BuUwtsfTCPfAm804abBBXS
jCfm2GwJGAYrNsAJUBHFRZoGUbMlB3T4+UiihP1rfbhyCNlAZbMvYtJF+1VEI38hl90LvNj0dMY6
4yntC0zPSoGBmAZwTM1z9tO/OVnJruCtR+URm/Xuf+aQf6UrUwkqUKLMymaf0caN+gKn3CDC/Nmq
ENioB3MtGnRAbEqFjUMuTcTBOEnQ/hSPjTdrOjupbEIe2zgYjR4ifkSLTKtxujKYaTpKTJbG+k+X
CVuRxtISEX4v0guEkhePuU+5zZnwJ1tuw63myar3zbGghxwzXPY2Rj+TVl5C9hz8FYsPLDkPnqJJ
GxwRc2QLwy1EWv+xQGhJfKFHpFKWGS2leR7zvbyikCKYuscnyLyFIR99saq0PcR+kLKVx6IVS6c1
O01lp0xEtVgi9CR/gx52COrXygJ05h9BimdNrwT3ii+M+rlHVNY6w1mUIxQIe16k+GCpOHP/nMxE
tLKvkTllFG6wIfma28bjy4SyJjJm4MXGYFtnsLH3EIRO81Owiz5vMcwKvElOMiZla5s5uTFCCXCa
bvRllH0TkWAWjovNN40bfEULPDJQ23sy9/G/98208+LyXPyU7oiFKH4ZVqwYJY5tUDGMsETYaeb3
qsYU796PiJMPbtJ2IFx3M2p/qU3OsAwllc3HGmW7VGGi0Hj+YgEUOFu/aCPmqy6ODyAPNc9pIRiX
aMsCBtOqCywGg8kytnx4/RQ+TUHnjmqkUwyVFVYq9xyf5agxL4Qd8v+PW8LmeVtgyOgoG0qnPKpl
KWD2AYR41TBRWkdSfpw843KTEs7Yk4H7UrTOPlbUqvnnWZ3nh5cX+L0xl9sMomP2n6+o+cWjg3Od
iyVCrCP4cxQ7UPwWrWCyzGdh9cPZTSAPooM7urxbWbpd37osivnT4bstI5fqy9DCRafjhv0xUq7b
kshmuGhiSGtwAdT4jSTheor9eSS4Mhoqsudx+u2AWBDUrZhmU3ynK37k5F2vqJgM/QJr2odNu+HD
hvDgYXtc0QMCPkENlJ+GPXoLhm+pkrqyls+R8a62MV0+uu2XjVIxnwjrPlV+AQCmr0D60qWXz/+H
vOcTJ74H77dgm8Ft7NxPtJQ7CS4dfg7IXm7Ab+1jOBY8+yhQ5YuP7zBGgEQjneMnLecOkyoLt9fS
i3/DvVWrrDNb0C876W/BnMM3CUerBG+u51/SINnFFklWZrUezUQjoOot2eQiSw7Uayi0sonl6tw9
9TN65teA3VOeBejWi4HrmYiKGxUHRkvTKAPY3wdgMp+wYsxdEhONr8G2AVS8yPgxsg3nfcdPiP89
/nVB4d+LIxO6lFganDfc5XU3xXJYJfhLVWMp+M6eRyxG8QU4Q6iilNjAzRZvu04UvQsSdCmTzDq2
azCs/LjVAxfU9m3rwFGqzMnLePkJiZz5zfEKIhXX1QzcXNPL2HShCT3HNM6kzJ32cNhqJbySrS0t
mvxQS/Ta3E5btKczXXKMOE24dWZB34tjA+szbtHNcuWxZbipKGdCdYigGNEsLxhVvL5yjLBmhrFG
zVkP9zQVmjvH4xLjgmX7oq5NHn+1Uiee4irNK+OKqUTxeKnKwP97tTOoesGlgzvT1CqaOl5n+cEB
/rBFVdEcm1uTHUUTL0mYCdBP15GyyzQQAaAExw2FcRPknpkrNFo2Ag6D8mrVXOgBZvnrxGtDatAm
YlgmppQNXwoPITmMkdPPGy/+BaswDoRsRn1oyT1mUv4ahU0y7a2B0yer+Ww/hAeqLGaJajrNh4Xx
+Xv2epf4BJPCiqy7VunrcsVg5z4LaUD6jr/yBtYl7cnMpBOJbUYkdyi1NWIx81CKeagHSqfquJYN
HHyQ5r2lQtT9ZpcUQh6a8A9bAebbqrulHfCK7Hdo0eM3hJTC2cTU1A0byCmqjnTejmiWNs/MnXKR
HX0/6TehvKVDB/5TYg3Dm2Zzyil8tZSQvyVViXh/Aj7AdQQqoKYbn5IEj9DM3ZZDc/TMuX2zdPXf
phjAdZk3IoQbjAM/TDtj2suPcMfFYiXea8FsQQxQ4HfrpwZcJXgAxDPe0MTkg/eK7FxEiSsQwv1x
FaSIwOuRl5DRZkHYcJ7j0TlemMXTAzftBAH9EKrpjqAsd1U0yvfrsuZDnZbYOJbOvuJ8B/zjtlMV
A3n6MqrnIbt5zF8TAIQ32gewXJ7CKXOqW7TNxtwoCT36qN6rHvtOSu4O+dqiK1vRQRqf9q5ocbbH
X2fZa6NgwH/iDeMkyPj2VKU92iRsHIRKWkVWDlLolkJu6a1C9L939DL55yK2nlnC1Dd0TtjLySN0
Z+/uIUfArfbo/bkvPq+AR8HA7FLFiPd2ns71KbXnqtTPK2WlZKbjaQJscymhN8CGYIzH16wnoES5
9D/LHbT/p90G6NdJI8C/jW150gEbJaY52xMwKnl7iq3PLbcP0RkYaixCpTjYn81s5rQhVHFelC0G
svmop5AqNSVp0eUbIgaMPsVDqDD3C9vNZeNLWNnZW3WCkARPjUwOfk8uJSWofUF4Nhj62fTrmyXs
lo/e4aLTpPrJ8nDgQZSAXXaxefgnSv93uLdsh9+4EP1nVioJxsFgyz6HKASoR7WgidpNbqDgBGEt
Uz7utgQwaaxSSScukSO7xBosLJvOdAsSj3DJT4fCFWImay6jzwMotfmmjQNA9YeZa3F6Q99KdXg/
wwNAM9NQzFHJ6Y9Y4cFMOvIrRdsn5AN5eC/vH9BHRxeIDzw1R+Ol5xFATSS1/cl5yXRRP+qS6wvj
Roe0LKrNdOilPQLr16zHW9eg/lhP1E/4+q5NwoDK+fuY9OqM23QZaWw3x9QZ3wHk+/KQzxYCsjr0
F8lvIV2dZxzIMc52O73p1piccg7ucL6uhmRSZAuzOAnZjaokVj20cLT2qPADhm1ICx8HQCCiIS4h
cUEh+1HV0p833WPvzEk7zyv70rMxB1WMoL7A+0EsWoA+N09xvx3+e7oUmlMuf4Aru5vJyp5mx0jl
dbRNvVSBf/6+ybRRUIfRhepjJXKZplOPBy8AEuEj3JK0NyVZRD3uQbMYnrFvxJKbqgL0eseEgYte
RGIMGad6+HasiQaQQzpaIOMuudvDsruSEEUk9MwHHOa5DAOwBzlKEsXMKWPJhiBu7tO2UCBkUEDw
AJ734+pnoGz8MACiTj2wLvf625ZtlWbteNk02y2UzGPhU/vrPZ184X9OS0Z3etyM6p10w0VwNAe3
+z4pF2xZjBDWGx2CQ1RjCxOUj/HCn55AML+rsP891nmPan5g0NGUyN37MxWqDdqFBsFBBFTNGkGj
PYy2bYNazS5YnIAGxQHoW+vShiC18q44TCrBrzqI+XZ39T020P/ajBLdtobo+E/jsVe03SzEVuOw
7g5Usg7m3Vq9AlSQBZZAjsb8UEuYUZMvT/QgQKzyUt7OLHMkZ4Efed14txPadQc9RYP2wt0vPFG+
+uzxbwm0XFzVkpOrx3tZlMMdsuKdAgJzNYJId0jWKujWH4Ajv5h3m4edCE1fYp54wfFPBJhwgxc9
LBhqzAMtiown+b9zrYEjQS7PEhgpWIafySQ/yQtYYxM/CWKC6aNmX/7iYXczkpEEnLumqP4xh7bm
Ip0GCmHz283mOQlxRiHmFvPt071KyNkEg6a+XXLV1I2DqtZ/wCrXyqUF5K+21mcitJaT8WNvCoQv
YJcL9AN9rT4K1u0N+wQi67ZSb/J41dhKmnJJ9hHRQOSymd8Nvk2v0pdBCs2FidVW8gEn0qdZk4CY
485OBJUdT77K3Ta/s3T6vDzZDde6RFZ7Vj4rcluf8WGlWMq8El4YEm/hqZ0pHBifIh/e8a6+QrAn
c4U16/IlCcjyXgNoZCZPol3tdfCybgPVB3osYwudrPw2DV5aVeRmLEaV39MkND3sIelpU3CLNsVJ
LbA5XC+0dYvStkuEaKFKsToB6rNNaBpSoP72OjzYOfm2S6uCfyEaGTC5HYFoqhF4EdWrD4YuoBN9
kp29CHtu417ox2Fz4vM4mezeqXGCZMwGjbx0WfyUn4wa8cvzbgaCY3sxlPdq9lSlg+uPqyDvfjQf
NOcXWi+IWGms8gyays66EDzXWARigVbNTjD8JizIcPx1ecvDPn/UQqKNV4Yvo5/eRdDsUCiadB+K
/5rG1bvc8M3Osnyii+Kjrma4fCc4o5OQp4NuWPbaEnfZ9rij1wFF5L6e0odYLkaKnTkQF5x/5y8z
+283hiJavGB//08cw2hW7e5bTToSmpBnZF3TqnuNjV6PPQD3e0TCUfa1ChSCtwmAZq7PBUWWx7HW
pl/BTzQSpncCLlnTy7jJ6Q9iUNLZgmidsJF31O35ENVa8vyrWQ7bNe5x8bF1gHUpeYxK7g/9u5bU
jp+ws6kmn0DkkJX8pusHCfJyzkaKBK8sdXJ8Jz2BkiSuFaxQNjaUjGiy7+EbPuB2foZgJLOE9ucA
niQRygWzKB4C4UQpTc7LvOFUT0werIo8hPrglFbKUmqWLlcAPs3VXbS/cChUZtf0C8b3+WsL2HTO
1JS6ev3dmhagmpfVQJesHZ2jhOHNkaomN4/K3aoHi7PWTZIqlx75O607YVdXcwrJD4ojD8wcGSB9
s6ef6zfYaWI8iflN6T0iCMpZidAeYBN3d/+lPjn/9KFeRjsLwzbZ5JtzsVGv9TOOIKFKTOi7K5Es
U8NFH4p0po7oSbHGTyr5zgyfoJfIwM9uHLGRli2ipr7Us1NSOhLYZYTJkg1dIzGLJwHFuIhLWW5h
VenPwdEQ3AkflfPhbK3TDyE8e2M4ZawOYYsr97oudKweoxQVezafCQEBZtldnZ1inxuNpp4chtrK
HR+G7Xaguj7MbNwylzT05Igi/E2xF/9vHDhOIHGPPLvSnowQF7gHlxqitZUtrgGqBdmLVdSEZwBx
RN+xFZIE9qjZfHSMZ5zlKCxzC3VgKtbg3qVCM2CtR9p4fS0nDHZUQUTVs0iF2gALqScgPUXImwPQ
8sbJuJGcrpG3RIdSbbt7WGTPsQkaZqngfOLse2+pnMsDExtPRSAqrgj6atzf0rccPld/qVlAI0ty
9HgSmBJj87L5RZiyp//nyU7muIlHRvLjORDuh9UUWZo2/v31eV7sxV2zAJDSZ2oMQaWxqpjU5L+y
STUxX/SaKwIMrQaTwyGFXsw3CnxivUvqL7PG5s5zNwuFFeufBpVhiGIk6258bosI7PuUakWlXmjG
lHIvYvoHyB4oJkqakMbeo05p3m686STJEpxsAiAN0nFEK3rqIqvpOMwW+f398ghN6Batm/Ygx8Eo
s2MIin7r0qBfYUTzXFPAZQPaFHwgJ7DdEWMAW+55/DS4ODJ5YNJJkt6s9JdQXn7Bj0/QbgjYsKNk
CHkW9d8p7/kA9J4NHYTRo16V9QLAsbmSwY+83HurAIudGF/sRgFsTBHbnnp3dSb5w2yvrN2a3M+T
D2/plZuiEZzmGuX7Is2AdpDOoIjHo2pVGPH3CUYYFJP8h5MG4uqFe/Up/R7h9Ozs+1kHxlZJ2LMh
5Ho25+bev8EFUWD2A2hOJUEqynMISxWcKVhHdtNo+hUhRpJxNoI5RmazgzHTG1wFMg8fvaRbd68o
mMtFq/X5Uo73G0qM8XdMx/jPy+/ZJEqdl7YfN82ir2GlrTTE9LSVkhBAUdzJXopR0CLamqKovy7B
Ipcjvkncau5ynfBBxOA427sRpmM5xDCwvW3BjVi8v3PhKPtpm82ro/U5a5g4thsnY/cd1EUbYVMJ
ZQAyC/xCUe+vIdWjkKvcAjVd+y51GPJYItnToE1gKJc+RTHse11tvB6Jlp8iKUb5PKqnxXF2Wnaw
UN0op6sSWdwDDS7uvzH+4GrvMLfzd/lSRfLEdY9PNDVaJnRLxdV7yg+L+Y7ZC2cINp9BeZMyYBCT
vNoFFIYHPei4wVCxeYzGoMXOI2PIwj+Y4QDbhoWPK5l2x4E1yLBtAA/p217Ne3AkgRVAA0wi7+dY
iYhs5gmHYPfmtfntjI2ruvQQy/TX+BjbbG/r2W5uTdpWDHSBNrp/oeRGfXEzh9hPy6aE95E+fVcT
MPRXZM9x4zO15f12AHTju0WzNDnWVHfCqOXfkxnV6bVCOxeM01+XnR4RChgLX5ZwFDFY98NfNHt3
0L1SAlXW4RpL29pBCmmXnIOPK+/URFKYkRJ4OD9x0c5i356JsCrZoMgJuXTDVvlNURPfAkeOPtpi
G3aVwHNzygss0QMPRBTFNy2O2y2KoSTH8GVz2rqfrmR5jcjvH7RrNuH35SuxwZKQfBmBEo/sGaTd
dGOk95MqAVrJPvFsLh2lAA0DSuRDUDohW5lmCo4kS8Da/Z6z8htW72LdH1NTDt35zatKa5nXxjv+
TIF0Ru+FiziyPiBbJa7uGTSwfAZk+kZ4ZG4GskAFC0YluGx5wHeoYtzThHRxeVEo5bugGYiv9c9H
DndZxyxnfEE6DxKNGkZMF+zMf7f6yczSw4UdthmRQh5e74qgpEOTSkV8WhUMPfBuVVNbeC1TtnWq
IAjNvbfNFZyWVDs8kDHwwX9yD9w5nTzF/PISm08Q8ehJR35Sd+/y6BRzJBigNTXpoGKP5hhCY9qC
1Bgxc8o9Gjl54M29Ce8I7fQJffFcEyKNWSkNioCFjySILC+tUMumQNE00Y6a12pl8urY3azM31WQ
5URWh7rA/qtghmxrZVdn/vRTLduiOn7YTBrE/Jw6UqrJph1jYlHnW/4GzURlwysVBrEunjnKzbfg
YdOOtQQOqya0e0XzkCMUYVR4vvaf74ayg6WjHMpAnONqKDrsSQcFhC/j+I1vx/Xx6xYqeZjoYhWv
c5uIWk9Gb33VoqSDaQALAlFUIj5fhaUYWkueZrnAaPcqZovIHeg3hAU5nfiA5nqkkxi4KBvfdNEW
4rHFoyKkVCL/bpAMaYbFgLrGMa9jYq97ii8pl3J8rcuQtUiOW9TWp5Ip9bDwf+gaIRDt91dgk7Zv
MkVNWRBZxsTOPiJ72tdNkcPy5m403Q7V3IlQAeA/I9cEelGm8YSbqkvkr6AWWfAoDTNptoB5dQBc
hm05P0Tc6OZoCpYqrmqiBwhInlKPlpbMDNJ8HE5gWtRxtei6rJLL98Ppfejb38kWlkLJ9OPGFjox
XXkbs4U3f0RH5C3S4t/1poBkaBw8Gc9sN34ba3E+sv3Bo9NpSRdV4HQUSIS4pecpIDnOfjTN14OP
9EJxq9vVvHl3L16L8ixkCOfvtjG9SUYS2RkBscoUsmiBp3088QFTpuz6Mhqv2yZpk9w+Xqx4u8F5
yXg3ldTXsskknHcOxj5sZ1lmAp+N003rsnEYpSXNUH8yDcW0djGDH6oxHhltoDeqXQPwGWjXruHT
MmYoq/s4yRgP8LWEBixGkMDErVzPJ5Nxkfwxj3N6LoRddikRl6jKfFz0PsUVbo+YlplbrzhmHBJQ
E8T2vycFeIPXNzF4F5qXMaAmaCl74K/sjrsMm2HhksYEkdygyb4NEq+prZ1a3YC5ODgJkZyBFOjf
VX/YW+Mg2RWiD19K8msVmFPoclJT1ndwMSTYrnzOpxcI5fKoBj45+ZH42t80Dv7naktgiJAmuFVy
qSb7s54BdXZQtaW1p/ZkDkL6C50ADOfE5XsW/AUl6sPlnTefaS5C5SxEw7VM1F4eUzg6FB5kJEAt
k//fKVsk77VOy9WqqG2afVFNxA8hFPXFiEMRQnVyA9eGkBvSQjr91KiV3IERMJHq8qtrV67DV33R
4wMgnEtL9Nc90q+PmcnxdKTT2CDA0ENHG+/LR7KrZb+3RamErHkdhmKQ5K7SlRZQwXN8cBBhWCRH
ErxwRhQ6SsSWwekgxWQcC6Kh06m6yfZbs+/Ryz1VcUxaDgLHy/renD2nbw4vC7yiiu8Mg5uDmj94
K2yOJs1n3ghiAr7VSYOr8HWunkea4G8B35xLhb852FSLVhB+ZKmCxsMLY8J/nsTSn02DHrAg5jlc
RGRUcMtDJIjiYmr/CeooEr3pJqAePktCluVdWQZTngYa4XqZX5KdVl4Ybzhi56gHM2EEbep9t1G/
l5H0L+jZ1RQBBIwU4FS+1nAOky5pmeVd30WtITLkc7Z+jfmk85Pl3+O3054NH/b8+h/OqWSuAfeP
m1d5q6gqjTZWU4zPQEstCgs7gnvsgFA9gPQ3OBLozvbThIqH/7N/MAwqaNOq4DAcuMWytYg5IWBu
c0NBjxVO78U+vMug8i8Yf6RNct9aVRxIPa88G49PoPDJiHamX/UXSDxWVaPuUAXlEORhXSNRaL87
JZ5meRMpIPQu3QyRT2XdDFx28H1vmkjN7iZUgQvmO1WOKsTw0LAtXUOIQsb0MavdG8mPUJfYK/ba
uPACkwlWdKgAsyvcvhi43wU5zzpOAvKVuY5DOLp3Qq790obdvUc9exTQMHrq6hn0y61pnGND2On8
6f9mu7wUTqlkLiU9jsYFEovdZHaWsUb4M7wXB+UylYbLDyOWJb3Ia/LDjnVhsfJagNYLXgmPiylz
k46G75Kw6Pm/QuIHDRUf8U4LBI8E88n3k2U8onXtKDvT7FlIJGUaDTWgJNrRVKyFnyaMLn+oZFp4
Z/N4tdOwPP3Ti4HCeGZVECz1L7gxXfBUh5cVXQVH2dNbLk3H9d7ZDqNdzBFp+XTIdHg0usiwQnPg
vWi+7W/x4UnEVB8r4ejd2ilG5Xy01uEQMb07R5SV9eW6a1JxTQWaCbozioE3HTAyYDRMTx3fd+hA
mCpOTK+EibzE8AOQ1woNITtM8UscMO+JH+j81cSrBhuD2ySQXTf//OYprFmPiV314YqIY1EBLKDE
JJqaITwOGrBsMJgKfI5fDhTB3K9mGobYdJ1lhPu69kFXiRXUJtZ0XInoEwkKn05gSzJZd174Yqjv
Mx+UL7HvXYwItCTYC6Kqdn24jtN6UlZMm2/zpfZ2XC9iz89ZqayxLcZBdphZY0EBFCYTmXzG2Ph9
01rIl1OLy/79glNTmNFLQqdvcHhMaolxQTNzD9B4Qc7CYrZjAmc9V+5vuZgUznCW+j8wY82vB5G1
I8PvjGiJLn+M5fw7+KrsxmsxnIDY6AZdGjIGpSjKVzYzJE6ayvDdrQAhzpzCtaXjQ4jCkMmGeO7H
Zi7eLkIkZEHYr2pktGKYEF2tAVg2/mUqGDoNyutg+xz45u+zs07vR/DBcoZQA5DPZ2rVmqYH/QYv
TXmPf9+D9tbP40G3MY7qAOYSHR6w+lDRgdOlE2GOpC8hxlHeQUpMHQxqKnH+gA3M0EEYMZ6xxFWT
PnmLeuIBzKhghvyVlP/1M2Nyg6iY+sdQbX7MslLXKue+gwo4swdCtv7YWCuUjBDhPLHGVUtprShj
XVyUlbFF5ZEAyZm4A3uLOBAD7fG3b2Qe/UxVy9BWZK1HodQWynqdimWlvwWNPaEDXuzkobmiLN8/
dh9zfSoqQouC62dF25W2XllRD0xc7T50HfQBcEJ13I2ObLJB+tWjMHDyVs3XhQWqknMrsJbfshcQ
XTfDGqF2e6JYX8sKvrALDS2JqThNWAENGBP/teZ2iYqm59GrYngNjckZ2JS2cgH0aCGNTrfZqOb4
qGARjTYDK/bKznu+wsi/o1u/TdkTvt9OPU+v3iMElBHZcgzWgvQ6VGlWLpSmV7vXMXJG8PgA/YpZ
ov9ZSaUuAjxFZUOj21zhmFuWFEbRJT6uKs/0Ybe22eiNUI4bUaR58Rz5D9PEgAXjw4foiL0+dvZ3
xkh8aYbrHaQRCGFcxAdYA4RH2gciI+aeQQHtUxx7Qe/mUxJIONXTSYrtUsH7HgkP3ZcwB17kqyG4
kENhSFXOagyz4qDsEfEklbEdRRytji2AObytWUbHflKfa9NnxBSrUBVxLdGRavup4k4EU+PyQ9O5
qQs21K6W8lQmWcrFRL9ZIzWfRzkvxgWzELvXFVOwsuBKhssO7fj09y089dXwwOlFpOVTU9JBOB2Q
JxfbI0ZHQUXQvuBGWP0XUdY73pFGKY7l897OzchxEGNYYIa1XwkaF6qjTjdx3H3ezIjKGAwLbxnJ
Uu9TW0SYC4kWr/+dkTx6X4bFvGlJAyc4KObsEoWmhMVMwywPNOfVY97mvq4/KFJEmSWvBRFmkyr9
GyPN6gWhRl0Y9HygGZzGqj9JLblcs1cKfSo6M5TiwjgZRhcm+eb0jS6dwMVvPEwHomNSxgggqDrk
8TcA0S6jP5kgZz5xM9jgtsinULZjOw0bztIAZ2/lYzEhOc7iLHUqZ+cfC/HXy8a+/yyI05FQat8p
LhZ+R+J58TP0RVvkDd/pzbQeMtaav1FWfdJ0HzCtpNHNo4ly9cBi7tdh/INPGirPPc9HpsxGyEX5
zEB5r7Q5S3G9+zEu1rLB5n1vBDGcyWR6dO04cAYcg0pTggy6m/Jl8FHGxuOG+sWc+EV9lLLhIixp
j3RBdzwn2F8BIN2YnQKKWa4RlPq/gQtfGFaDEx7BT0SxxybLEZP+RAGs5J37PXyfmJe59pQ41GmP
7IKYqeIi9AtvJ+UEQar8YQFFpXeNoND3Jiri+khcmv5oAKtqvFbuhCbY512giQ9NfvF5N7ab6fiJ
rYec+9lL7iID9ZkVeMxvzmoKowqR1KwQPVCBM+jJhoQlo6lecIBE2X3U15bVXfuHWzGm5yjq8fqw
2VFI6EtYSFKxwnlUUJNaYeZBants85Lym7UkkyQHJv+2Ax/owFSsSYd94VBbdRS9TFMyCaaxpSGd
h4hpIyo3TlFIWIsWv0QPFa4Mwik52n3pJ7EpNUrTxdvYwNWusPzL03QjJo9bnyfwl/KTP6Q8wsQz
ffo7uyYUkxq5LtrUkzjcPTRC9DkC2/IMfzqC3mm47JVTaro8alESp03OAoEZm2R5hDmkdMex/arn
Y5uvaKAqn52Vc6raDZ0RfSW1+lKo7ie/gPAUbAowT9Y26nCQ7f6A2pt8NCdCFSQaxRWjFXjy8QZi
TbdfVbSzdlk9MD9wA8jMx03XGp8foIU9Yq1kU8BOUeM3p3knHpUKDFLWgFYBlGIx/AHvMsYoEz7q
SfFiYvaoGlyi77Od4wZZqjY1doy0uvlR/vin5KFgcSqnTv/RhBmXQr1Ro8uYSNPPSA+fSRtUZO81
oPv4sD1bYeiwAjHk5jkdk++5V6GbDYXRJuopASuJ658emlQcaq/CHDf836fQGpECVyz4WddzDPCJ
GfPkndVl2kOF7hEl56bZsHgNjD8IFzZjeBLrzKlvCCRrwyznY8nQVklskx7tAHEAgKjEQG65UWeQ
J2PKfwWX/mkz8K/+MMwbTwBOa6sLhahdR91xlnR5DnvXt6j3bn7C+n6CQAfQxuD5LAPkqKmdFz3a
wVfEHZPiHCzEflUf923QsVFS+2i3m9gummp2e+A84/QzdLRQpqZ85GUTFDv+K9D74/yVobZy9Mu9
KmcsUY5xwuWimdOOtJVcN++8M2wiP6zHZ3iCPFY8Vo3H2A35opzZrtThcZ1pqyRFyEycyfXLcSD0
aRv3ZCB9rEnhujdg6PjOASmw8jjVwjE5Tl7CzkX5CAk6pgX13TfDZXbxZEBfjH9ijI6JJcQ5nMjE
b1wHLf97zUD1dD9dQ1dGhnkMinvwb8YwcKZFBsDW1U5WNSt0HrMfn8v5dhlj1pCP0nRaEsj6PASf
9HP33jOVnM5aNpYmb1z/UhnPsMri8l5+k4TXBLwANdCNoncuHHy948Qt4xKoGTBH2s8noqoSWTXk
gAN/TOkqsEPhTEUuInSnayOOWEtzeNMnSQh/u4+6hnb0uaiD3hytVB7gcbu/U8gctL5n8cuN+P9F
F3SYzpi9sZ7aYGUODmEYWtIQc83TFjqrZEzqxF7JGWwXkWN9yWFBhbHfV9BQ0VtcH8smi0ke1gzs
JSDqHF/ixck5ZPREw9IrRyCW40QRjlORJJToh1MW64v661b5bnAMPJwkY2QhYD/3hZJDUSpLKalB
e/Uyt8tSUxiTwUDzf46NOrKdtZengaRhtnjGHG4fZxLTX4/caFJdWyesLMs0w7oEV7FKvq7zpIs5
WnNDuonSDPQkyK1Jt3JLevPxDbVSZ0qenOX+7thug9KiFKYIdKqGXTzkcTHUN6KtHCSPEyXVTkso
VedqRECSX7C0BxVyaWejOIgyJKExjyoGZ69tBTayOior4BHu9aYbDj/CSR6aSvnWmfFnNfpcfdpi
JSkt4rLNG2tXtrcZL5jtVF8Ycjo+8yn4UU1YfHAhOfL+vcXi65EK/fnnU6TbD3AgW4K+4vVNhtwx
065Y5k9ciEhNmwWFl15RC3VBIDNNmSnxLk8ScGautn5MwNVZSAn79ii97+COhhzNNij4oI7dc9dO
CRGSnsqoEOUzUOAoGVIUwbOmZ4JYdt25aOOk/7cVCMksEuhon5HZh+ImO+lqjChuSUqKSDCboNQ8
iN4qnuFT5VGi/7Yh8p1cu35VWsUvLsQ3jIU57sp2JeKmF1BNWGf5/dj4y/QjPjvnyNxWqjXyfzvj
8oStgLzWRma33pn6aviIGDGknnyjBQY5JzazEPk0uZSuOLvFTlIG4mgUI5YDlUfiuZ9QFXTNl8YJ
AZyZgEbEUA9scf0pVdyaGX4D8L7uEpgdmoMu7mBAjC418CdwZYE54dXx7LtiaTGpqfleF6MWimAg
8z7uErDgtaxlTDGjt6PvFdjfGHs/XPh66aXPLjUaTJppaUG8Ge6ZuhKIlBatJMr6Oo2+BfCRMIR4
fKdi3qFVOUabMF5sZQNevotOIeVxbf8sPStjOMCQxAroXE69J8s/AcISS0Y4HhqF+4eRIR2iQ32T
gjzpLiO1vOgqGLt/8rMlLL5tBHmC91OCnnCQAHhWao5x1Tq0bxJZFxs56TJ20Do4WQ5GPTQP29DP
Mo1x2c1mCSLVZMNzj0YKKyzeAfiJH3lmWYLAqCZ7rK5pTJWoNC09lQmb9yup3DZ3mIvHY4Sx7v5b
azwK3bUvNYMIIaAcwscjSh2/cTzMAe/dNKRMIe8/JQMlGmtj23U8mVHAMN6wwsZefD07G41JEEqV
ep/vf+iEusMaWl/qgJa+VANHCCaQilbVQo97VhmCSX/An98wusnaZCJUnEFZcJZvEqCGXyiLaRD0
8ac1nZNLCZy09WG9lVGsH9NaZ929R0gac9sWATziimj7dd4aeypCxtcAMQEgNCeIiPDhBcamaAWz
OOhUkeB0Bpi3MUlfkAI+WmyHOAVBGZpLnBGm7G9I0r+3axTp/Quxoluhu7kmgGL7G7LZ+cQgZGPR
Y0hnuRMbdLXo6tcVChEAgzn8xunNIq4cgeZeNTEQWlA7yEnhpIuiCeIaf410pX2Blx6LWgNGyhI0
DZUb9wtFJHdI+E+cI7ZrQ/P3crNf7zkkzxT/tgpMIzszYIwHwCS9RvB2XO8RfRWAbeBgWkNRkga3
TNJm9fiRj5tr4WsQ1y5WbwQAUwoVbxXJko8pfGlmq9oSop/zCfx+O0o5o226zA3Z+SBTVLCZHJDf
epW7USyvoUKQuTy3kmtgA42Fxl37FFg4sMMHmU0EHBz3NVLMo/QQBzzEnz74rOe/IncvHCgMg9i1
X8VROFkcmfng5qb8Yn1rZn+gSNPKcZLl7hrVzzU2nuZagZNxdDOb1c4VlX9aKs+iFCyprJe5ghRq
ukR8yK9zrw6mCGX03b99cHtNCjxkxG1g/AJnBPrcsly2X6XX9mkrZ9LuzXZrKMkcgAvNprU1FClU
V/bbhznwTzdc9PiZguK9rL2sc3EGHTQwE/SraNnjRExVwwpPNteCA029jiI3hXEGApTntGPA4WUA
H0Z610q+OeCfvCuE1BFXnXhhVIsqvKHIB+dsSzIMb/HrPBbFEbhZyun4ukU3oHeNNWLlyF5QL2ro
13KeEi/Tu5vQil6KdJFSOZmGQZLR55QqY5WckvBTDWpjcshKTtYn1e6t0/sDm5bMFRFvAFFj+WxP
vWYztSc3I+uB1nPzd2eqnNRvkpC1VXCcIyTO17OjV0+0GCMMSF5R0jC+YYq0ch+GCRNlk0qfcC5L
6McUEBGSkQ5A6WWIYTEfd1DCM60Yju82Ap3BBFC2jL79ll3hJe60tSBMIJJVk61wOOAl0Osm9Z+p
u0UwUcxweA1UOUIrylcZrre0ydlicysqfuR2HvOEe32rtzC15r3BoR0s9vhWj/sby1Y4PxJ1siGc
RWVWdJtgm0NFcCshkfLz2mI79rUo/AKnpFCvoyhLSWeWzhjnt0f6aefsRWMlCp1GVEitmP5zELs8
iRTy4VeQwItF+erdmy5kCBtRzsbZ3bT3DJweZhZJnsmkcbC26xAk/BDrkYLNbDNsi9aJkKi3y937
fSEis5NdUlNWU3dzrQkOiBMDoPSlydvDf+f3fg4W9rNhA3djBjr5gPuhOAHJTOnNVdgNJ63gEfGR
Nji+5tjESra3fuyB23irODMwb1bAdEv8Wgs+ZhRaOZVThevNB2K3bEx+tTtM3QfMUFDgUHJI7Q5c
9kjSt4A9/cuFNFhmzJ4eBa7ThRmL90bs3cpUlt370ncQRrqkX+sl8XO6+p5sKYGv8imy5ixz4Fx0
5Mf+5b4KXyhRHcRM7nMCkTO+quwvWUZn0mreUWNK2aBNR3tFtnQcjFNE8oYPpIk0Lt+2l9wYPlIh
HoaNHhfpmMegJ1siohwOrBFjg078CdCjrCJjw0Jnzc13y4dCgB3Z0peHqbM2hvYkqDQw5ZHGdwu6
Jrx8VR8kqGfyJusEv47MzBRuHppkhRM1pesPPb07vPoxnZK3425nfRVsEo2Klm5JSHtAbG1VOiyl
6ukUgzXEOhgZl1yJgjKHHGNf5csf49VgPQx2h4g7wv/SuINIA5Omn7iihkpFou0qiXMqOmjIkRGX
kkvkIZFjA6NxLYRlmYpHh1iDFc1Kmic6XjRfDFbEF0iuwpgsKG+PoBOrsR7Br8O2ITpHl4VjIpgg
uLV1CPfGHb9duNk3YB51WQ5hZsnagf1I1LaUV6BJuwZV8Rgg/iVN3pcwd2Iw4jgDWcd66mKzytqw
Y8rPl9R7aUHkunypiF4NSYGck109BdB+CIur/1NSrI5qavyS8hrZ8IuGtbpsYKBrV+Rhiu5OVdja
Aag2YZq28vXeYTfFmDe54/yzRwkU7sFHUQZGGEbPoGaF4laFUob5q5g9mL3opZ5o3rMB7q80ayOw
VWzPj2ryrO7Kerc2LA+gAbkB7pCxbvS6ZlC+O4IXHYbTbET3L3VPagDidk2Y3iPv/LAJzS+XiS8r
GJv1HliVrcJVHmVOXS0DQZA8eRf4ix1JRgOmGfgq7JSJbHIQvTytkM7Q1Mt3q0EPH+Zvy0j2Fdw4
jOP1DqhqQuYsBZSqDa1TdUgSHJx+JfXdYDIdKrTubaCUkXCYxfD+XO4sUdmBm87N3sjz7ZImMJG+
88XjuDpSRN5T/IrRvP/frn4zWxKPhQZyLrlCuCXvWwSSl0ZAhls0Y5hLrwat5KReIekg+mcMGMeg
eTqjVJN8o+c8RSlTk9BP/bYJAf/vkio+IskECghwfA4p7HaOXTT8p3CvsdXg6wbjNPxG+JxsyMXb
j5CDOvSyEzVSQecQVoMfsvFk3eq/VvIf0aI4i73g28qRtCXZuijxRSf/0wMiWq0HEh5gxxZbWrHI
/quBxHml1oFTXGh0w1vseYKAgvzlYqIv0nEd4/Y98THd/tOvMxJDf1taCQWoE43rEjrZSQtIMm4N
gwwYDMNa9koI/ytgH6+9TH+st5MPKYfXlbutFSHzwbMqGQ38WpqznNy/l3RJn2EqO6nq3+zsqXha
TPAPLBiC8vcie7dg1rwqe2I5M1AqyeUiqKl6XKrpmTJkU4JV+4SXY2zicwxqmG168JpuAnFLOHCC
lALgtW5MGsYEbi4YCeQJqtysKA9nJJKznD55agDCVMpqVKHFMh1vWUd2kirb9xGWlJh8Ql+t7QX8
A+Jj+2yzOGIMQe4YY48uv5dFSCmOOQOF2jvaMlZZEYP5EuWFVbiVfPiM9AJ7JPBKVHZ2nb+6R0eQ
avNYl56eSpEsh9W4XFobIw6LdkZNx2XZ8WkjQvY0wLu9/Gcf9uG3k3/zLf2PP9rOOOsg3UVr0jxD
tjPfG26yuqSuPOBbNJwgeZxcPN45tn91BS686zOG5rlYFWvCA28BREmPo+cHJ7XhxUC31CW6JjKG
4X8xeUY8ydGWSblFNjRLjlfXkMMkfj6NfDBDchaDNMHfIAcDYEcFDLiD3L9hRZ5HHhl36eiml4FE
vUJFpZyVPyGwkm+ac0Sbb4AV/vsZOBj5dvlXryQty/TKl0He336r5ub6jcEGZh/ikDWGMiucgRal
GUqPt+i1i5bmjLziMOUZh6FjB76LRERYs77ZFVXHRmgNoMY9UNH4z3fnH4Eypp7dKgDFMNu5cQZk
GMT3ST0wokA/rtHKS4ExfKt0GbnY5pWOS7oZSMulgpiZKnkBn2MtgFcCRqqKF6j9rGdXaTYXSkqA
cH5e21ESmA4GI8056gZuvNSb96FFvkdW91MsS3K7p+oUE7NwMuts9amHsBWs+kSEh7bRT51t2pPL
T7N9O3N7HXGePQdvFPB4+Z8smYPMs0F9jjsMhqkp1mDWUyy+xLdO+MxIiBHfs5IZaY9qIz8myzFM
KGqbOs2pewWXkSB3wkR6qQLIe1CYGz91owazWYZdJmBlWf1SCIsHLEBsPPTEM0Lrn9W/9UyJq5+o
Hw6nIU3otgMY7687S2/FVD9OIwMpK/Yn1HrhsCfwPOV05peRuFRqZ8keKbyjTGVKlvIpvUB+9YoC
JBKEmfaqblO6nEUtcek2kaqVzkbKbncjxQA2GHbweUbG4IqeVSWHkW/SziuA0FOsqkEO2eBqQvO0
kY6fT2czveQczsKYhikvRRC70MfUJYSej+9EAW8PTAqNJuo46dfmkTVsqrVPPIh/tMWQdVIq2m1j
gZ7IPY8QmKNcNBRkt9ropckkWfaECtvi6zikpLMvZsrP8SGe4yQMOjF95Pn+lKnJdZE6WvP1OJ2S
Bd+MtvK8nZ7yZtx4tHNeTuUApyerDFipFzXvWi5vXRy/aMqHvBEjoZ7DKXzoHuapZjDTGCJpR4Xd
ddMN8mcbdnzIdeQyLCR7K3f0RI0dAhq7X6D73OeXYZCZWyNRlD55eWeZqr9iiDlRg2AkYz72i/HP
U6jNbgLcL7RoyRo1RTf9/zx8ojzrpovg4jBsJumfXncnIUwA2+RVoFhG6arW0B7Dmi59wc9X9Xjl
Me5vg97pkxQc1OsRx9UrUi4TCQkWxIVzfwxxzn6Zh0JAxbm9Tb3DCVamrEJ2dwrRTy5QlR29+62K
/BT7sSngg0JIDPXdWnS5XGUz/2yaUTTlCTPfBZs180vrjOYvxKH0tTVblWzPOOjtrhmlgN+WmN4+
xtw8AiQ11hytv46whxvB0kzI+wYf+rh8R2vPxzbj4xMViUHPIsDuUbzDKQxvmecPbkVJC8t2A5vZ
OmrROdBFqd5woupLs11NGGozrx8jW8HQBeUY5cMF0fKqqGqmuF99RyxpnCMbJ0bKi/8esjm1KRpT
759nRiPe/Xd1y2I5+u+DimzJR0Ml/Kg/29N0pQojhdAYcNgmxYA/CllgfIQuu3RYdq11nKUeUgW7
pxMNrkMIWavijNPhQASNslzTo3tWOK33vZh50mTXq+ys6N7Mq4MKl3WMwwbo/4UcEq1cs1eCNY+b
tq0Cl2FZH6+YaWlXwZ8OJ307OVMZe5xYRWEdRu0LYD32Rr4fvKsgrkfkttYL8PxosguPJf8j6GTc
Utq8GJLqTO0TMWFyhq+V9WfCU/tJ7bO2NsivjSupu3nVeNYz08hITq/49EqpwxCoztMhyBOoYk0T
UGPHWGOME0FFEEbTK+Z+W2JIXdlOf5I4OwMmMO7uTCJVaqqgPWD/KZoI/+/+fZCI6MOqCO7TfuWH
JjRHyuSMkRxsaLgr6nezQae+Y6BMALjicb4GVJdrLCCbVrAknKhhaYRK8dHSk5na+HYFn9BaQx5q
iuhoPXm/kCOvYwj922Sz2gqDDH0tGVpS+ONxps+lXmIqmAo0PWmcR1q3LJ3ISq1ljyv5fV/pA9Po
XnZ/LTgnZrfx7fPGRzatgh63DH+sTcYoGah+4AQOTUOs3+mWAebCe7a8zGiCGvYUHG9IwGzyAYCU
L31v+2aj6Vo1rjz7EPZ2oNvHAVO8N+3peXaa2DlqL8swN2YMlgJ5X29TYkdJtiGTTTdAwyVqX74u
jURZSwEng2DnGojiSFK4Fkbd3scECV7mf8Mdp9PK0e/K7vyC3FDhlysWLZxCKIEMzMHdYX9e6R+2
QPkEeAvOXORMM/VKJLCw0AQAOqIVSDxGCZNuyUOjZoYET485UPdAXLUBcUU2h+vhnE6X/eLK2Sze
Z/dakT4icY877zd3N72Tx43WfyYZ6Bd8y495xbBJfXdT46wYamXfCpJGFVyTs2cNR83i1whXD3Vj
atnqaTlwS9Tz+4WgT5QydbGIXELSs+pU8IUs3ppyiMtiH+tKdN8IAMGV9li/g+ddRKhs4If/6NfY
lsn6Y3+iN7pvjogXxslVACqrIo0lnbWQO9TOapydKJnyQN1c2Qpwurtdxj0UVS+tbrrihKx8bhBx
sOLmJIp82hUsEJj6/xqnO3oVw4j1v2XZRzSeEhcVSyAGar1gEpXVOt8wzbr0Jj6xFMTvhVM0jrb4
UAXdwaN55WXqlvwueSqNkH6UAqSuqrPqIwcmimEOXjRPwKOLpbqG6FLpI6YpBknG44wRR/cxpZ+u
/+zNkNj6I2+YAxltpVbuQEYDPkavf16VT6PwkTnwHPT7v3lV29FccQc/H6ck9rubfJ3iqDenvssv
SHoYddf00nwr2xspd/vAFx/v4Q8hqDBZVsSklh17rjBVdrCXipRY87Ac9wv5WUxj2OliXgXg3p02
nTHgMZgKypIbiJAFUKgjcUxyrMwUda9F7WgCktL+xN5fmQhnVm57s2xpj556/JAYuQcwK7ceUOJ5
apr4vlm20YUXGbYw2guDNKc812GMqF94PkTH4Lc4W0WMCcJpvRga3M4pFyNnZy0fxIUkE8+Pwxwi
94fi2DmFCudX76Rqjaaj8XlbOc6sx2OWpRRopHJywwWVSzh3Ry8z3unhQqzXm/jp8sFuUPraTt7F
m3obFX66aDdPClDiQJEsL9xY/WUlmnOdRRs18OuBFVCnfSYTJ3b7RzDL1VRpvAV/6r4yRiew2vHB
qQaIoeG991TVfUGWWTP8LPYkHp1xwc32g2DQbcXR/zOzbydagoUWrdfC//J8pSGFiOw6HU3hSlMf
2tpvi27h0BOjw/Zl8JWsINk4zkIgT0D4nbHa4G7bc74RadjBQXIwu+bQ/UrlropDfbrUCXnX5tqi
g5mK5PEzn2KsNjUF6XQ0nOKr6DoDj42bngZ3/G6jEq6rrqozjm2LUGNzz1D7C4o5dxAq1cKaOIek
Hjblwr2uayCeNJ/eJFqw88KT7UeRDIHuBo1k9WyJzLVcYv29beqSDcPk0StC3HalcznZJWnqJKcN
LeOa0S3TZ6o0yuj5Po2JU4pPRmfuTdVZtoGrQweYLr9PJvaufNdeHzpUY2JfQQS5ihFmOg0AYC2/
qkw8HHf3Gla/h5FtseMTMskXTjkDEvKPlHDL11Apk6oT4A+YdKlkjeP8chL1RWfEMce0KQQELisL
bU2O66ML6nuN4JJpmUc8ZVlDtPsJmg0bd+jwAU/fuagjTlf/LSSYzqRmSt4ibsqmL5JHvXSeDK77
6h1F/btE12RNPeZkhWGezsgfzco9fhJX2oUS9hz2AamIUUEJx1dSlsRG8AkVEB/J0LzChi71dsIr
PlTx8Zlr7lkJF3kJm19pfSE3WVmdwYYqlPrfv1MKbfkcDpN9mzYNin0Q5dP1tqtyxoyqmuxJNDfk
xNGsEPPXuymMEbRt15HzwtwpMvNkXXBzm909d4tVMcJwYCsCdW0xivkW5FPJX7Du+fM5vjEMQjOV
n+SvL4vJ49ke0Q4AeKPgUl/NzJXkhH+Na/eKLrJcr+dNT1qRF+3F5yanTfVaYWDKwU0W3B4VpMGw
J4yDFrSf0YTg1HdIZ28c7u3a6xNvxYEvLAuVVvWBYv/6g0lGvKZmAk4Eyqi4fOiWNqPo5pELlYjR
VZrROHbV9FhYcm6ppKQsMLjLNB4DdxWaz7vNFWXqZC+ds3ceuvfHQfJ6chGHaX9OWeHwUD1ugOfd
3qKpu8QaJ6VxiNnFWRi6nqp/iXQXZoszmifgU17fjFr9P+2SxlRhyLlsWq4CWuUi3RhDt21cwD+6
4f5gE4ocyBR88qZ6lU1UIXbbwXFSzzV7ozI+fCtiUUsiyjvkeClOV2vJJt92dPe6aX11nGPLhej0
LrS/ZMDDCUpZJ0qUmiJAFsUKCUxCNvNy3VPRkBOinsjnoILKM89TEkUpA78K53JINZ+0Letq1Ygm
5vr52td3fujBQRK4Afjr6uPjQn1HRX24b+Le8XSIITq3PUdxhCgFxuIxalWH5VDqhGYmBh5kV9J1
nwmA0BPoN5F28rNmTOCMjffsC+eDCRNpfZVaTLtEacFjQ/g+fi4nZPxibQ54fQbeCBrg9BHuC3Ll
kQsYzOyxItWubKcA+YgcUEJgnu410rbwKvE9XM5Ipxt2w3Kik9paDf0M4ICNjhf/Kta9RtJufZml
rcwahUIy+dm/6CWiMErwiiJ/+Xsj3gIxodTdyRa6MCWnQREiSSyYbIFQXHTS6y+Qvh1KJeglXn0o
o9ueH55JA+nQj4PqXgNU4TnWJiFrsNbE777ujLnUFrV+hiHfctfgoWgY0rqiWp0UK3tmRP+sVSfF
bUZMlOKHmOPxhoYm2PUlrJHJ7InKSCTGS370ac1CM7rOm9swg7sJdAQGuOPm7ZicTwLVamuqZH+Y
C3Me8wUeTra80QKyzRqRxVuzfR4rkPSX3zpeEkaFwdnbuJjaEhY/olYKp5UjzNsnNh5YgecZPx7K
lVN4PgF73JNEMkZ4jrS+/q0THbfEhEv0v/5bUb8y9Xo0tVRildJixA1pj3A0/qXgqEwepCzBx2dx
UKZrbRfkkgITY1aTxMNv43nZ0Rwxupd6APVnZVRP/dzUhA7jSeXcUM/JPPospC5rP8FSc8KOxCMC
vppn/4hQMSKRD7VGt2dR1nxNOdS25BnQ2Mr8kOwaNiWvjpY4WMHekuYFmgODKztgp0kxwNb4w+Qi
kIaAN3BDLPDgt7ck5J7zDA4OC5D1DcjgEIYdCcKnLoWmytSYBRNv9gzxoCEJVXUTPDd+eheuRLDT
8G59l0H9Z81CGPA64p1/lm29dj5E8cNsLiVUv4x3faISZhGt7Qr5TSv+3RczMMYyimqvrar6AJ+P
uBacfCTYSPA5OYdrURJtkiHkLkxWGasKpobezbmeCEUb4ZAAb4Ygxmqk9SEAfNH01jBEtQn3xsE3
FOrhY61ykkZ+c3BY7tPaEUMyME1j1BHpr5OuoVGRcCHNC0xwiYeg32/V/hfUT8wATunWgGzNXfYZ
A5tt2qBGiGrisG14l3pZ4QplGF4/SZGbl7G/uKH7f+PZt+PvhH8guQHz0v9f6KnSpRJpHAfDbgIY
MzRD9dq8+va2nwOxmCdgt0RuPgKbK6F0bKlFZwQfUB170O0t1C1sA4Iuv0qQaW7kJUXJqIcdNE7H
xQtSqOJDCKqkehC2hxtaDdYQby0fN/edJZkkLKTEFPlPIG3NyIUTy0ZE5nxXmBgjQzw4NinlRE9y
qlq4hgA+gvm1rYxGBpy2E/IfAe4EZg76UrzFUDzzoB+pu77WRhtcjaOVg1c1D1tJJbZOORABDPxR
lleZe1Epit5DJHJ54Sw1kUSvSlDizcrvRnvJrmKNn6uVzPsqDiCYLcEJQdwAI+Dk1XR4Vh98BCKc
tspnz7LFMwO8XLhumMyQRplAMU8nQE776cdbS5wfVAzSyGvQ8w/TcCRrIa72nBt7CWIn1GuIzR5K
fOXPaJj+brZ/EIi7ZFyxrONK3e1rjuG+BO7NUfqImGN0ltEbLcP+1T304pObXSVFRdvfqPI+Rrdz
HFwPeZLaP0YRsFmTxqu2XdKaBPkD1qQekgxzvAsoNJY7DIPTe1+Y2eerX+A4gv3uLawd+qlfg41H
c8RS01vwruviMlVNqHhSJ5zA6xw8cwRzhjs1kkVipQnHJQWTiK9oZ04FR3o4t55Bp0paGjBRpneY
Hb2frfhYCo4JkxsTg66D8rraXkyNmeO4E3rlYtGja6C3W39b88Me2PtHUcUdQ2U6xaO6ve6d+b/x
5HcmKvnlMQp9jUMO3dQ9AwJj3Tca+ru4oG8sP2dIrJyW02VL0Q+qDI5h/cOI0elbr8S5/71HA4tW
wyloH+PlImQGjA6FkB51QQ7ca7cH5eXqP+YsqYgPMnhV8iIQEUaDu6NYV0p5KQ3+llBIo+Oda879
t4XkbVCHKgtcwxOoLaYThIJEt/ycCbwKi3xdCv7N5V7UOlpX7arazTvI/M3x/kWfHXtRUmMHPYJ1
7Hd7UtATKzY2jZZeNccgh0xkT52HTrrUrK8QeTAmsPBTSz1Rv90HB0IKdq7KU1p3APhStYPpKkYl
FKw2r1zn6ArFds7JtrEDk7STaFRel1Un8KpQJR8iEQ9FC9gA0XDW0nX7elgc/CA8PCmIcbedsE0l
jL+oM4Y6ZwSBR6YD2mEhjqJ/8TWDRuHNA4Y+CtP4QLsigmrxSlqNIYDPuOblUsl9nkPwmIIlmcxw
QqPcZKyky66PB9F9DyZF049wO6xAyXVdPo9V62K+DjCBbA4cBm67ZmM1wLazyv4pgWjUKTaGE5Ip
/UU6NO+XerxcVRSUayF1/Iu7cp8ho5AwCXEQ9f+82+obx8bGy9UnVjNFHhfy7ta1T6P7vD7uMbv4
Qm7sMTngNdiwbz5/hzPvTxXz2LpK11oT63pwwjcJ+Y4VVV3s5u4UNv0HHggfUz1ldBldQoC3N+EC
j5935fBO5Zo/4cC9XJ9Djlnd8KMP4kDwDZFMzn4xlui2VcNWSa8f8YFl14Ljwd68bFxI2F9yuk52
zSqzQ6sHZ+SqkhjfY+mxY0ua+G2j5PiMOeWsxIKssZlLHrvmq01npEFIPOrpqHu4OlD0CHRtfR7K
BnLTlWERoC+IRB0BYyKlfzfalD3ZGPjFXzF6MnL4vfxrLvmVJdRrVc8fMq5J+4kVSSxixbN1Nh6z
7gB1bV76EFGSaRFFIMtK5/eEwNByiNbzBtFoOmkQGFw0IWLWWO/CErWWmBSLldHOrx4sUhN3SoNo
jHwYJCj1XfcRFaoSIziVskc7u0DFZJds/LrkLeiyFL9QVRv6Bz5udiOiq2rNCIrBrZbfYj+vfzPE
RUYgRSlkHbvV81TMXByI59NWTMBb1d3Rqze8kVl5Cdr9R9OcH3KyCMvGGCx71L2093nKEcskJn7K
iFeSqq+4eWGDh3DsjvMHmnL+yK2EMiqebaC416l2aIRK9nU05Ik5BE4wc3KVrXVK3/U4C578yZjX
Z8GXFLQZzoqh4XeSF9yZdBBmO/oVkgBnkv9jnFey7PSD2orZrQBXneLLM1mChh249vLMjLjX+8Dx
GDy0PBzCZvWzUdANUUv2ImsG8JqZxVqYkKZkrZx+59VrbYBUTrmU0+selJGAQv7GCsa2ADp6ohSn
8peMKPnWZexEX6lnEEIi5X6x3OWB2YR2RrGd3yozZwMMNOKDa9QWg2ZngaqbYQ/IjFxBHd24OAon
wCcn3V3Rad6iWcBc3Mzn+xhgxick0UB0N4LOMuBlfZTZyt8DwSFnSw8tDWylpMZQefX6Xk4+a1pv
EkYzSzBuLyabWkJTG2cvGof5kstkwfMqWiIwAleROKwRp8w7JAb05w1zx15G7dLiZJtNOdDyXNNv
TM+V/YmHOSJ5++pSkLaZx3G9ALkcVkzcnjZQu9ao3BGPdoAv/jqVBBP0Ngnb+/AQ64hElMlQ5pDS
vE9GVjNC5ZDluIQ6qjKhMg3iXpsBIAOYuwCjWCFkHED07R+JyLZS3MaVJZ3Ck1lnayJDv/jLtp/f
Kro4utyMxKD5S5b8iwoVMcZBf2FAvndmmEliUjAN+8yqUFu3mCK6lSaWsBAXu0EloTZV0lRBdtJS
la0g6N1sKmkPdejRUhSsDg5nUl/9USTKCpTeVHZ13iOK8TloNQXAinTvjKH3iRiWLFCAIjASzg7r
kV+sGALPVdRxX9vyrgvAeukdOWkjbLjHGULXdMr7XjVVOV6RxT1kH3fP31oISuyIxrsapeKzsS77
h9nOWYWyUrd2fjXiefdtNvJmQoHjJmmvey31pHFdEP+fNTGGmghZM7MZ3821Nt1R9UsLONavS1Eu
Vs0YAEVFyf8Y7KB66KvXzkU4u2swD2kduo6L2WFJEMukAvBVDZolwinG3KpZ0BNNXdoLPUzFaL2r
lQW0XeIeyBu0AZAU6A/tkyG29Fn1fbGFFJJu6SvYl4WEANqOdpG9unCD0zQgEmaz3l51y4gYn+TU
6vQjUj0XmMvx5nIrjlck7Z4/6wKESEqFvgmyKXa2DszYHjV43Uft4LSf7HwUYT7qd1x6d9EMJNfn
Zf0cOakuaMZcxRyQil60a95yrujNvkTr5qZo1F7GKFev7OEFPp4hCe5ztLw+Zkee1h+JQBhUkxNB
a7AuQtV8kGko3Nj+O5vU98jHehl1BLUVu76wEvUz57UD/fnVfHkNfh6TKr4Y6LXR352fQ3Hk1OBj
ET8TAJy5HbIf5SqyvZ1fV8m8FORcNbFJYr7Lxd75Td6GdFTUpHIT7LTFRZ3BwlWndIjkh9/KvgmF
luGbEUgWtjPypNo/WKom7C9o3PTA4oh5Ycky7F8nQK53iKIL1mA30TeIDs8Pc8fBsXizx2mq0hUF
7IBeC9rlDX4Oo5pwYlQHXB2MT4GeuwJD27g/YyerecAxgMFrT0VSet0IETCuuDomuIuWWa7LCM4q
tVzyjjirBkPBPwxdqeYqB7AfK2irX5B4Eb4FDMHPOsAQhpru35YM95JQHlj8i6I5/PVVNI0Yv63d
kgQtRN+OZ2NpFrePBmpG1OYsJYS//ZMkwbCoo4iKJxFM14brY6N1l1BCqfV27Xuaj/wG2ueJy86P
J+sA7vqTG0N8hKXEcgA8O8piMQg/0An2AkYD11apaGXYEbUFBTY1/lfK3ZHdx6haIsM9IrdDESu2
IJLRu7//DDWRs3Qy2cSsjEKj7pewytqVRxD/ephaJVKeJwfeV9InJgwuB6Sgx09r9OnnT+fyZRtu
2ZBUxa4Nb3ChTKvZOoVW/LoYrzRi/1k0SExQi9P6kWkt6VrJfHCG7wtfTHBemEs5vW5uNlmCuEP5
voAzRLc7El/cb7NzAYUWv8wiI26x262ffkuk18UNQdrR6HPpjt2ekLTKEdSjD09zKAC8KtFTCjBt
uNcIAlBwAdYmlUcPBhfwBdPbRY4wwlK/COq5FyIv+Fpsm0Z02PpkgB2qrZcj6OLeilHyhJqV+7Yd
9TGRAKbaHksqJV6+WEzguS69lyw99E/eHaOJmcOGADMSeBhuOAJLv2JHiZZYlffFzPirLjs/1qRA
lE4zyUMOaqftY+pwWhilJxtREhdh95T2C0KMfdNWi+TpJLRojMDgi47W3fXwG1L0af4sWKtIUd9o
7Gtor83v6BpvU8nUQca5TSWabw+FFJ67evM8QAnGGFrTxLi4W/ye28kgCEMFlMJypZ9J/C8XA+Ot
vMySsBbvHfjXly3/Z1JE8e67pe3aYMm/XYvP3s8PJSRyeq5e+obJCwOu8z+0bPlZBjWpjjXSJ9ba
8mU2PW1yhNZhNYl1Y2iLqqqOhhTySjYiXbzBemDzpasd8kkhHeaoV5hhoX64B0QGVDcRccyu4Yd7
sBMAlFRecmKG1HnMJ2VZ8ue8ya7hbXIVA3GNn4Ws/Hv8pz5mRb0tw3YkAIgp4mRWVHpqAltchFlk
Ipc745bolxxyRgx3JcCI0stAKOl4DKAQ0/FJaGM7dERUO2ETxUIG1wSmWcRnkLfGVYrYq7eTWDmB
N4zT4BiCVjjdaKPm4X3CLpfT6OCR0/Ffr4IOVQO4a9LMNa9ybRLN8ArJhKrDPCF5UheW3wdPey1B
iuUM80gUhm+BhOUqUdnF8d0tDh4xYncP67cst6aQNZ1WJdrioR4T6V25ktOBzs9i2zGo97YXua79
rO7aZH3o3YAlBWm6dbbL81wGouGuN4ajONKhT3h1on4YoQV2hW1vAM0WUgYZG78g+TX6KMWqTxgq
CbutUaDCr2E50Dgmyum/Ep1g7v5Qzs4h58iQ9Z/eg8aGHu6YCHkWOwyBRwrnITzYzMMeK32vQGIB
8z4bJ1z4dBKGfjibfL0qjUyy+/4DEUYn9zRR4aZfe125E7+rCREE1C32xJQvQGfYFulPYgFej+dS
e1oRSi+GGL+a5J3w1wabexbbG3mjWOH/uvp2UloAvz6b6JtrJnkVQZVSHUzs4f1+Y0L2KBm1YAr9
pS4QcqWrT0bllu630ou7YL+Rp1cHeSc2mbmaV3HaeruhczdDT0tPvq1mzIz3L1FKVbDq85X9FOIt
cnSY+0tlS4htSXMV9lW4kMsgYZbY1GVlG4jqJy5v8fixYHrLIoyis6kPLuoL1b9mSV60Zt3Yi1q4
kElwTrd7cB1P++MXTRzWYcvfJ/B+kchBa+FVT1jTX0pZG3nahATV7t6RCRVxpCzkyuOQhIIT+AZF
0XmS4tVBThDKcPybohaYac4SaykjIZnYX0DfU3+n5Tif/pb+IF6yi8BjEmlTuQpjMh8w7Vm+0AvB
irnMApHuwWFHfgjFJM1imZ5ftgUDquRKgMOmwo0BVoq4op5R909S/i9ck9PTVUBpVhB21bgn6S9n
rjw8wPb849qt8PLOw0gBiE2c1XIaI82tG2rYUzzUSSg1I5hRvCwF7kkCY1XaDqi5GSB93GAouhwy
DBPICq3pUTNgwNb96K/TMDTpFBjb0Bvn3qyXVnzob00lc4F0HTQJvzflWjsRumI+u58bCUxk6c2A
HfDT8g1qgqrBXVmGvsDT55A2sOp8Y5F/Hi3onMMdGyNQRP5jkxL9uvEckwJ8O9wM385x/w+rt10N
c9zZTwA+70NwnhBcB2dF/nvrWLMbk0sd6Z4HNuLo6MD7mZu3wTFTi6lU75EBKuqcUEHTHRBRVjbr
k+cssh5YF2PYc7ZZLdW2MHhFkaqAMnLLLhS9NCx1bMqHZJXdwf2GnsbV/sU7okrZ/PgQqtxv3szG
ivdXAYfVMeRMvOVwohm5Juk2QOdQZR25vJ7HdCLljMNpFPwBzmCSoI2Lvnt9oH1EPCzbWcCFpaD/
leRbo7+Nzx4FYjqMXatj38hXlzlHFeMKeGXvjnAC+2873YCI7HodedDpUUzfcQ8Gcv1SBVv0O9su
G0nqD85OUIftGWPS/0bekJR7X5ZGFSQAQR4qZr4xeAqiFnmIsExVHQoD54eTvvvQ7Q0AWCADK7EQ
PQAf+O1dzO2I/e0vCzwCesluHlVh7MPWff7JWxaosiV9P2H9dcMzXfM7T+1pg13WaSPUUckn/F45
MPspqCHDoEUi0npmXW/fA8LZHYc8BoH22f2ByuMtwHkhuhLSSEYPbkUnk5wKoczCD1QuCuj1gmoo
8ZokUV9JhIWNFN4GBd7wf9WPCxvWM5z421Sd6V2pJI1VnwABM4z+GO+yoDTGUpPHhTDAG3jvXKjo
q0zihQbKByxxL7b2FrAFAafB4mdZdP3fKwppQBU8qlmm9CrjQTJhKxZErHOG3MvN5u/UuDYYoNSP
8i1Q/QxtH+9nlDEeQNQvkrwCSw6ks7rcs98kaMyZBeT5vkmjv9bGs/bCWjGWNU/+EoIg7oM68nKZ
3bE6LmItsG+n405vEATEtk/kcZKdlNPwHzTEDrqyT8ixWcsrnFxQY5vb6Lu51+ORIRumdEs2yo4T
IpbCFx3VU7zeaWIGEK+rf0qqNnmIHHXZ9SXp4cR365iYJDNXnYD1XM6S8ECSLyqxl8EBcFvi96qY
AztDC4vDE9A4cQ0jzdavE6hMewABJ95qEfXyJh4idCvf4pmjVuD4dMMwmjoA/cD/SBQ4ml7N4YB3
qjBF9b3v8xeGL2IqDL1zSpEqmINld5RxUkZQ/5UfgfXbJ3QY/Kifxa/J974W/+xbHMk8qaw9abKz
UiQhG2d+gApoAxsJ80U4S5Rj6W4Wftz23vh3yqAfYVDj4g/tusPcZSpyNs7m8eGstjrgSgVGd9nH
zxAevnKMmgL0aJEoCd1D44ZBCesHe7itm4nq9ZDKfDYCKSctxGwyu+qqn6ax+GKm8d2Z6TJOJi/u
Zk4dth4vX+nUnh4MSzQqLtBM0LzJA31O1PMBpTdxW9kStlF98vPPG/UBDUgO8yfKEoRBrl3ISows
dTSlvb3ZbVcJk4hcu+zsY4F6m+t94l5eUsZo7ACeuPjxYzW3Lxs6RFPdK08pIjPCHRINPrkN2IXw
FM2MMFnWDuD2wBNS3Hrc98EtsvhY03TpSbzYBOoyJTNmHldpy2fXDNF/xrMpjbuh7f8nFDzBHkZF
jfarQOIy2o75L6axWVeu/Dm79L+tlOT3kgi8SwXzoJOB6SADNEKPMaQq2cxm4R8wn/T+PINzJP/J
H5nVJ1boja3LHUDfCIEbzItp+aA5xXqutNZrHDuq+3d8PIP9uY1FSaNZr/rgwY+zamVJsDaPQK6F
O4PlZcb67fhq74z2Q2gZvC2rjH34lEKEzTAbnf1d+lvGs42ln/F6PMbJhInfuva3VgiIgb/kVvqS
UFETdKi4v8ruLWSfqh8NRhiYhf0SEIdqKwEDCoVGAsqZyECykCnutJRVcHJIk0VPoNMSmtRZ8RRO
nV86fruOTEBdax7ExEgx/qBxXN4AS5HzNl/klrTnh+L3iDwHOJg30TAa/hCnod0FRAQFmQgVMqny
jo6MkCFdVVC34wTiDh+yV/ZJmbN4O0HNV7KeGNZG2yqABuuTrq4DuRut1YB4NerB5XMeLdj9FZ93
CXC0aJMi7n8IThFWX4c/vgY4xy+5nW6EvbMVg9sE+yc25EOLCfoRPz4YEGt14ADrl9EfToOFlqzU
Fs/3iB6RH9YDo72Ff878SJXhlM4lCFjjJGtaXt6qNiC8pYnmNjHiqD7cBID+mJTfA3n9AcEhk5+V
ct3gjLeMmgygr3w3xsfBr4Bzn0GDJMPmFtECYavW66ea6G//JKuPdBIEI0EuIXz+hlVJDsu8NzlD
cOBLVZR1hi4cOGdzUcrhsYLmFdviqoZOdthmdJBHh9tzarVQprHqGKHsdSbOP60TElQRHZBvVEmS
aHl5rFgjouM2EWeLdn4S733UTR9M28/PSL+WVrJOGoo8X1alLO/egNbYtQhKO6l7r8aBTTL4njPa
D+UikMQgUcrQGtdkdEtfU1fsxY2VgbXYYk32lEZfmETDsM9PEMS5PNlPJgAaTRWc72pkWU8IcP/l
3ZoV54muQZCPSfSJGALy/xeVYkZRPNEJGJNU+gitUTP3dNEi9Z65Qu9hhrXE9k8VqWqT0zJfvKg5
ov4n8NFMdOIFktCHzpBwfwFNGociiiKGMaV6XW1/1pvFUoDhecdJuvqegLDm0T9KScUyTSOREjyA
fLl8APO6Bao2UQ7WfuDfbOOS9gvii4gKtiriT6Yjb7xBC7xQCgLQ8E5WGb6Pxr8LbVN47x1uslax
45eIEtqkpPICwpCYgILMISTPbIwvoFEvNtUF62J1QtOPOp9ulMBChpTf+lF+KNFyFUaa6t8/+/Yw
6gGfIVnX1+yTL2jIRsSd8uuMpJ2/t5170yqS7pATt/RU4RHW6nVg6ZLanUjxt996qKVZQovRJsP6
PR5TDiWjKCLqAdM6nDnNF9reHlrfd5iKf16Oy7Ro2u4z81oAhfl9kHSfagQ6bytMCsdvJe6v+5vj
pqvhCb+ONd1awH0y3flKyhqSd83jyCeHUTqH9X118v+p6x0kxeRzhW20j7jqNm60YhjGdDo/7cWT
Zzojx1Q4kEb08lqC8Yp9XKymDzIdNcpHqfzlwDtlpEF9S2Mtll7/TdW5broFB+9stCpK0ASk4OvR
yFM1ocIyAk4oIPIo5irXoBvI1MVGFRDXfJgXkueYLu1iLgKkENelJqmA/aGTsFxAsIrrMmtVimxj
aXq9fbQX1/Jni+84nuo6v/xB5kG4kAols5HvU7klV/j+zMrnovOo7ZM25YJYXH16+BS+Ntof6ptM
hCruEBgQNoeakRUScr5v2ktMKbi/bklZfMbHij3iEMBOLnx3ipN6h8jJpnRupy87LIyxlpyOBQ/b
Om7GaIHgnV7VhLLfVXWhF8Ze5Dsrsjal4nBMzY1oeM2Ws3jx00+bUSogJb4HM6OSEqGZER+/su+8
qGigRZovG44TXrlRI6WWMdlf+PYE8HD4aiAXuH6xIL53SzmUvebVaO6d2V8Lc4mt4kYBkemteJy8
vosAlwOs/rLJKf+hFuF4lAdy28PoPdNSKxqA+pUIEwnktrU3IT0vNfo7x/d/QPOKsRx900xkyP1I
EEY6lHu3WqLA5uc07cdD2i7tKZ/6p5NTlmE7qEdPRpEIncBO4q414agZk1MNr5pDe4/xSBzDnLG8
Ezn9niv0o5iKnMzSaX2yUx7c/jkWyhJF20pd5i3xQmhkTsab0f8/Uq7se82jRX/NOyLjOmL4p7Bs
w1PrmJwkaxAdQGwMOgPTdhQejL922obuHvIdRsogyQjLeK6hBcWW3rgz6q01shKJZk4aIn65fkJr
IBI8Na18CSqoL5ceITQ26ixO6VE+mr8oZ0H5sd9NNDmTqcUIoz6pbWVIKUNDkMTaR/69o+TFLatp
Yh0e99J7S2kBw1j4p3TpoJp6r942Sw4d1RQrljYAAu4Thnz/4DGme7C8rAktSvJFQGihG3UnXosu
WCuCT/OB+8JHRsmqsS9ddFvLeOa/P5CE7tR2ZvbjDzLH4gaPVV1ELF+je3mAYXdlQSttjwsjqXFA
ULtYXriYzqLVIZEK39Lw4tehvsw8ZAnNiguUynjYbC2KO9MIT4+yLOuiHhC2v+jWiVaJdjOOEJEv
VzuuGrtzRNM85mo32PfhRhkmzB0zzSm1XQFYw14uSV8r1MFbKEfK7YeCGeXNcNjGuaxWm85MMVi0
nKWYRQS7miw5UJwJZ1Cl9bCxf6IZxMLjbeOumLKKHMnJgxznI98SUJ70omya6qO4i2j5dpNotr+p
jt8EWfX5cXkyxWhZs3rX7F6/9/rP6DWDMzAZ91SuNBoHGXvFhd94q+rAddy3z7oKyuGXbqtDnStK
3VTjh5YLm+xNzo7n7E1koXszzb5LTJeciMuUWjb++x9sCFHtxw0qA1qsvKUDdEYU5JqnRv/OCez/
LirpjT1unZxfHSFCGX2IDucd85Z8AilpyYOvsHMN6A7bwd3eiVUnRGC+iMgLMD6CGIRKX2/e4Abx
iWI3+JMH9loSOYM9P92FGyM+J5Hw+4PAXyg5KzgC3CfHH29ehSAKZUKfE9JQfbhukBCyK/dAHhUK
7tReIeVDFas8Y/U2hmM8MWWZli7apG32l7h+f/K0aKjXzhgHAr01QK3a8y/j1eppdTHm7j7co8kC
NDOvCMmZpY0cTRehXQxwY1Cs4MDPcLRafWgTnP3RIEGZoMVp2e8DEyvIg9mCvTpf15K0ZOFGco+E
Mob9AvoWm4WDlOs0yw8ewlpjMrM4B6pC+dma8kIk/OR54ZjSnN8KqX7Kd0KmqeNxNZfRRIN57D2E
vuuyrAddR0G+KM5FDj2gK6WdAq8oHrEy2jnaSoqSKHvA9qCzxCo4dfThx8tcrNE+uo298BHhbNV/
xUGz4A3lqVXrep0A1Hd9tjXMpVi/KqCyYaKvnmIolu/OETd5SzKfTdG5z8Ls6lycNz1odI/h05XA
wmREh3YVR3OKmE/HvH/dXHVvIXnaVgOepy67Oc4znt9p8qpLF/E0GuSdupfd1025qL5wrfv6L1lI
p4VOQ6jUFo8KZRjgdfkT6SNPJUu3JG6en8NxR3VsMxL7MUWAdB3d9d+ba+UZt8QOiYvxh8qwB5HO
/reDPl18n1dCrXAPkCw1LotlaYsQecwZX4ENCjbJmNTMyMBIm+MmczzzbtqB1m1B+gPXiCfsiN5P
DMt3mbs8x7zn5yAvpgXEWIRxJB95xIE9fAJDYiUzSocqFSCa9aDtiZ8OgmPCv6VM5o6db/sl2Dk3
Ri3p8H7S5djLh/L0mtS0lCSqcSCUSOx7Pb1iVnacjD7CsjXea40B2k695+2CQwqry7e+T1OmLzwQ
5I5QUFrK3uSVvyUagG8QG55JMwC1aTVT89Y7jGfmH96nQUhxqnUFONWigeBgaT598brfqcCqKoyC
qhn+E0O7e8WatONV7UEh4VeUDrejX/G8UM1lK/BvkSh2udyr0AG7nMQS/kcEkSO5M4AB8sAtGJ03
Jp2Coei2zRfmXMvwBm1GIsAQom8/a1WYH0AzwxBHyBwcOfzXZB/t8jfHCrfMhu5vwyKIuNsXTt/Y
bBVaYhOUEB1seNCJWNoWDByR4WkPjMQAlApGIPf9jF9kXBJ1LvYkceBu8LCLIXc+bz9z6Dr//7Tg
jsxZa7vSUa1dVvdE1Gxszglf6cjP3X4UW2KwCyITzEy1Va8NmwmMBgzwRxesvHzATX9IzrZM3pbk
/p++0EWRKmTAULyfmUbNj1sLzVVmJ8AH5RXXmDoSmIUECMQDs62F4zcmSI9I5+ARx4Cyrhti//de
HObLgI7NNnzO7Kfy9T8dZMt/OUi3jViw4ccPx6mcBtuOhHFFSidrr7iVeghOr/N4lodF7nsyFE+4
WtYyxPi3uXYnsf3STllZDs420lzF7PfPQk5nuLG+o9qxwU3ruofm1mLa6ybS+PA+f+T7uLIFJ7aE
9wryBfuXOibbkf09tO3vptMa7rT7TZGlVtBJllUl0s5f8n4Nxh0F5jx6CGJXWsk+XTNkRxw6scY/
lNlh8KvAjeY9iQwZsAhgTe0Yd7iNY6ecMUA0++02RyDyX9LZv1CxvvuGhiY2a+mUoR4bWr01lz75
o2s5nRTGDVtJVvvsscVF7j2mR6zgLl2td0/DpDu09u1w3Wb1XHh3gh+Oqh0R+B3U2ZcUKfLhpP+x
xNz9pAdr2Nz7nwTsnEY3Bpqdw1IjTvwzhFblYi6IaxYLTgpqdLjwsKFfDYy3qGq376edug99k0FR
BtJQFOlOohfFHSsYUutUKBoBI/LY7lEPZ90A/ShWfYsj21L8pk3bwlo4d5z2ZQjsbE6XYYdFLVeL
AV4Z1RQYNT9jvGqlwT/Gvj9K4L6uby6yozbEFNTVcRW4Upf2qur6l3+RPrPdGlUfOfRfmY1L2XEZ
yE+avSeIuvx51rDV6ka2oFAbT1xx6xrv5drCTvfKb+yuca5VnYipOXnPjCSf05HJWbPGtHQauWxN
RxGfpkAPXJgEC1qk/VI4J2doLTE+f2ZpOI/Nj/x29u0gvU3TDAplR/PN/5hz/gfgXITvreawTq6w
asp0DRz5uIuOnPazT4uWNA0SsVzQJtB5SwE/TnasaIl6p1eEw1PQV/p4E7VQTZ4Za22D+aCEUP9V
MCx2r56NBxJcSQAia5yzbj/Ilk1N/bnfz/pkb3XZcujlNU5EXB6axD7kk9XjnQvVvJgB33oRp8kN
uKkJQ+hjJzliH/X0CaRHkJhsGuembcF0qdC2e6Dr1mHcAUJSr6VCnNBu+9j8n5tPZG0YFpWqpvnX
EhDTNxrlMFMG0HNBUnO3F+saKEQwGkCmaP04f52CRagPiboY2MrniEmEnQlfO0IzJErdn5D66CEv
YuYdLtYvCuwVajQPc5cJ6kNHGw4Nn3bwsKYxG/0MW6bRi2VKQpCgZClKLDRcySRUh09Fo2k2dtO8
YPb2N4FLLY8TzvL357zLHoOZnoPeE4r2vv37lXwPn7ik5tQeTDr21gXHkc76I/WL4yI0Wm5g4srG
V8BRxLvGOYMKG5G44p5Ty2Wx1yQYqLmgeZujvoNXxePp3CqfTvZ+T1r3IycjZWGCGDKwgHcO2hnq
cWo/ElPcTQ/Gn/tjRmJAONDyw8XwXBeSsqLQcRJq0vn+ryBPH5FEpIO054kl8vQlGEdNceWtmffA
e4geK1HK7OzKqxJpmMH8AlyYxUNAhqmXXA+vp/dLann+AaRhYWnQbt57CT0exfoCpEEhFXXGNp4O
v9cedWozuaAMHjeC/SlFgeK1jzZVC+3q3k3p55+5fU07WvR9MiHw6NpP7BFmTFjSEvg5r78poJB6
cvjkyLhqJ/CyjZt1GlFz4wFs0bVfH4tq/L1o8y3VLy+PxXRyiTKyNCSuvM48rmgOHowH5eq4csFP
jouYcTrlefOAZGWIK3xiteMQIIxnE4HxHTMcQED5SMyvFIhyADiNX35qeZgB2njIXiyXQoutNr/v
Ietb6SZSYIryu/KSk3eGTCgf87PauyuzeTXDUSSlq0+kU7GPXEJ9biMHg1Nmh1lI7QKICKQVzAtS
yTGQMeSg4FcV0ca6587l72CXyLwsdedjeg2/BZqnWnaNRwPTLjx1STVfMTg4lj2mcoBpJL2ED1qu
hK8a0NWbc+btfbv9/hktME4A3r4ztl+kOurzGVWk4V5pxbK4hTcHhPLRowXylP5dHGDvcOjqNbhl
+aesaljoh7G618eUhOdTYRKc9xhqxFZbrnUQGfHiLuBl2ZsLpPpSfEfQKTV8q8+F2GMZkavn34Ou
aWqmtPjK+b9eFuqdYFzWRZfM3w1Mg6iloC1k2t0i8B3oIBKKKuUJhSbnFHa05uuOxrH5xtLPIxC/
YRVh1OngPgzKrl/AFvWnq7c/5EhGcDa/EaVnYckAK/V/9I+Is52ovptZDTsiazwC8IOyzuWXMQSp
t9XhB0jN6MsZ/XjyJN84CAYCyjuA9aEBggPPdy8xw2ffEUsXTeYeX5yzMK49bjegUqOWqNB5ty0z
u+GqkQkYxU6xslnRLVLUQXG/oKXalHfEiSkXfCzHKxd2fAVk0XnsczDlCXfJ+PywcRbdVVMzjQ2J
ArXUky1wf7Br0KdX6bc7G/kzLt42f9Zq9LBiCewTiOPiwS5t3QPoG+DKhMe+NSw4Kk2zqQoheQ/6
G/9q1LiGIDpYQBD/S+1pVKGuFhk9PN5QNMgZtMTfUB1P9SV9U+SXu55pgWXzjysyni+sJW8OSVC5
rlFEJ0y/9tC3BWNABZmpHwawBgH6fWNbkZt1PaMl+UJuULkPRMervX7WkTENpj4qGmky2lsBlFp2
iK5TJl+BgPhcqj0GWe0x2CRRYaDDQGmBYA3lsFwdFU9V0uxmsaXLPnpveKVdAgw1r2ms5SQF3war
hUiJkNG//+dTfCSpVI2DiIm9FLhghFR8Euktp3lXwYtzPS9n6gsCjqSrmd69TtSC6lnKmvi2Dgxy
zKMS53Kp8Bma9tFgwnkxKKkl1uPV+uASigrPNznsrI3QoF72VZ7CchJmpxVEDRLIJfyll4kZhSuH
xzdvwzxEzG75uEc+c3Z0Puf+IjEGelbnVo1I1wbY/rFm6avy8CGAm5Fd1ySdat3RtFQneav1bdQX
6ei/eEyhd176nc7FENhOsRFNFspc21slv7T4wY7yiW5AmR4ubQ5j/OW7ZcLfFf1nEDszyC2di0zX
CtGwdtGUIQgiWapZJhTvaphMS2glhkVCorE3VRHDlujMoX2qqyT3253WFt8UZlhMVMm5OCqzGRCT
AhLZwVHnLYjM+iaIrOa6NWvM+RK4ErGqaDqjLRln8okS4wOzzjygUjTQKi81CFej1Lkz7BtMBOvS
3mFtWqRIWH5cZLcNARB68vV/MCUxbt11e9v92l3Qm03bqzM6daj+JouSi1VM50EWE+LEx7/5a1t9
TMCfxLWDo3VjpCOhWEUN/s5bM1oNmw2+8m6w6AJ4dS3o2lgo5PPpwQF2VHy+9qwgzNegaiIuyexe
l2FfpqJdKPZ+dZxgtwfTRHO47TkYaEci9QUTeWm30rQeopzFzgaTXhW1yupIQ9Px+xp+6eD37MI3
W19cWFaWJKsa8u5P0kb/BiGWbPK/vqVVZiRt8dvpdeB41PlRr45kLy1BdjTWbNKfefctS8Bfjw6P
/ngpq11b+itmyatwmrq4z0LET1ldPEmbu7QiFjupiXOA1mTvaltdwhfsgO+haxSlVBzPtbUkNsDJ
bIf3b5q1w1rqX2NoyXH2xBmJ1wXNUbtmBoRh800rKIJD3zYv/mNtliJgWI7RKCWEEugCZ5wG0em9
FHE9xhwt0XCVH6I8wNxcIYvBNDP1cspIVWcaylbBoZQ4XtdFw4ymyeZO2QXr/KkflP6Udbx9wnj5
U3HB+EBa6M4IhY2pSAX9geN5uv+2YuwU9GdUd1YMnVVu7fqbmcaWKsj2YKE3ykDRhckkGw6vMJRx
BSDhPB+pPzilVOLP/AUnpysWtL5cBJfqsE6G74VMtPL6NiDgh7qvk+AxyseGnFRpCsWex5a6Oqh+
0besf8M6Yv4si+SJY/LIPaYovzZ4iOUu/rp68V2saSLOhNRSv4A5U0cuie2jBs/urJ9HqXXLki9R
yy43nEP0MOVtcQOHhmRokJdK8uZLu3s6EhPXBHwDe5x5UNGw6Y8E1wbMT8i2fdGs9IjXYt/KgUf6
PbNUroIVKcRctvCQfENw1yG07ZNp45qzq395eDC/LDbMD2HjvYPKXACp2d/a38l9fe3rz+FxcAZB
O99XOHUrl9LJnEGeJXCk/SPbujPY/PVqzIBpwrLkLV0N/E4cIQ4nHHnI9mNdEPKUHUIZBi+PLY5i
aHFqKE/DJ91HTR0TxPryhlQsJJwhzs+aaYdaElEbHaWAu3WTNl+9jHSfY19EiFXeiSjJAo5nhSHq
CuKfkIv2j9UgsJLpWm/ar5DqH2vggWZ6oDy50UGSYlC9VESkuX7nIqLES/5Q99HJCfRbCtbWPcMa
IEqt2cUYL2hH14hWXi/ai4hjjbuNmra2k7OhO87MdE6cb90fZFfFIDj/IAYjoOSkrqqiZNkNlAqN
L3xd04gTsCZ8IxnsuKDueRX1NIWN6T5yqCJn2XZMmY4v/XCf/01W9/65e79nJudxz5OLX9DaYeAW
wBaRpNvOf7tl2z+UKGtH3EDLNP+JFRDLvRamcV9UNiB4gtkvmSYs8OtRcUH9fuVEIINiaI0wYpfb
Xw6M3J/OleJ9CSkVsV81iF8H5WXYnCG4MATJXEMNa4zriAHJS2dgI443px5RWyeaHGNDT0fTlVhp
w6e7jHYV5LnEICKT9y5fNm9fuzZJ3kRvMHvEl91NlMQKMPG/dc366bjfMbFHHGxKi3fge/t/oil5
u6mGdzvwXfIAw7+CnkBayicC5XdqNU4Myobhpt8Mii6z37vbJydlMZBYvOZzQf1O93S4lMwk5PmS
MenY+hVzQzL2hZGG8p13ux4ofPPUK8DSd+KvgIQ1VdHOSK98T9v+gXOrxgI3EuGgyhgYF1UqFvvV
/Evg23/W4vv7r20yVAeQql5jof4Ku6I1S4HRc7eVkjE3/xpdNlRDjzljCfCOwKTfzZEdxH5Q2fHJ
tPNnZKF9xnXIkxCPbZRV7Jev+DDHRmdnaHIKG7r9+0E5ZVwxaVv1ulHbas8gGG3b4Tcw4ecZys51
/41y24izqO1rAH0UJ4yLkB/4rJCFO2MTAq3d6kSf1Gk3Wo3NTeaaekP8jfc0xNvvmltHtkgTmtwJ
sW1XS0XgRxMcLhfdD+w/1LGcXpzTCXct06bFM8D2vNHqeDyWYwRSs/8IQYCNNwJ10aAJBPmwg5qt
Dq27igjsT9MsWRzMFIVHBmsRJ6ElP6ayBwXIglF1HfmPaz0OX8a22wt2dcLB5W1xW45mb3Fl2OV6
OLS6MZt7BKP7RVbAjb7upWNW8v1xfN6LAhwO/zXhyOAjT+TFLeFggI69pYiYb9HKjO+qDYAXk2Q8
7jBTvuQiA8Vml8yHbS/bNvVpZfAzcof92+7dt0ufG/hjlJ8ygOmTQEiF82yIg0leBkJIq6zttF0u
Ty6uLQNIA5hZj87vxVUjKbLQ/huJBLow+az11TIvjGjwfO5bmq7DkTvudGZFRwXjw3Se33L+jhPI
e2Xkz6Bh3zQh5MrFiaJisSJq4GpyDBfx/MLTWKZY9x6oQyM4wk011UzNINdns3c7MwvJs1yrwP6R
IeIk5vwkzlyZmCqav//vK9AMqp6Y9E0Sl5kKZObm7JsNJqQXdJsPMqT/dcVusVOY0Dme/ukCW4pN
eQfAEnSlTJXkwK81cR4N/eQQUJMzAeOLwCO91DR5gHqg6XFPrJb+D13VkHbYHJ6c4kwDCGSfDsHF
369WfOn9s0pGDJ6gtqkwTINzLjT79MKqdQ2H6fgm5cYO3vTW2yb7wvQH2W55WABOGgJJH9T7KdeN
3Jp196oWfXevov7a7JrY+42Yie3ysD3MKWkOcruzWwIf5JcrndIdYqY8BVgvcJKkaZjW+tfpPhno
HpgHJcbQF9ihz5pHaPemSYMSC69eBE/Jx8qNvnoRGn6fIXPW1g1ZTPQtk1hvW7S6z07Kdb2qEcfx
sPFFKfIhaQPnFZkQi5n+JFbu99YcUTSbhv1BvVkM02Q/imfJmtvf/wXlw93OMfuAy5gL/BfNapIY
YjGYdJywKEfBALEOT8CP0dOo5t/emMx5FCJtBZC07dCgoLT7ykISgtoan/zESTwbp4x9SJI52M8Q
vfZQPYzvuDDQ+Srn29NYiTTbv4g4h6gR6CRJWzcY2X3tBxcdy6Fe/eskCosacZ7NfXbjOtF8CF1h
CkDoWtZB0FiGLojXWhq1MyXcQN7Zb8ImqUpN793BWMbEsCk32izPb1Nr0G8HmmKuujMam12tfPda
HjkNWgc9ohNo8CGVDdOh9nJhq2XdBsB+4Leu+US/H7Lm6yBNIxjC0bInn8bu0JZIeQXAPHjBlUpp
kSsDYCR4yo0NgY50r+egIhuaTmvcOblIqbMzthnpNdKqxb3JQcgoW8wrHu/cYQPNDvLUKQucL2+f
hLWmScx5C6HxUu9cO9Io3j8N9UImJlnhxZhaepdiQ6XYVwalsZ7D+Z3Sxpjjri0H07FL2F0evC7N
SU0y/NffOB8ZARwqFisAV3+xE/89yNSg993YvfzmkQ7vpuZm9lebCPS6Wuefsby7RPQXr6tscgio
PSs9OuSIYN9BoI/raoM43sLMmOJvF145JisvhNQQh5lhQo4cV9ZQnzjErW9nbO88/oveBI/X6GI9
wFmy5RuHV1rr7px2HeNYWNI2ZBDn+Adn/5+WzUzKOhcEs0CRCL/A+5jfsb+J7gZmO5DLPHaW2aAE
FtPP0f/LOJt0em7W6DbC5b5Pw/ktjSFVno97Iu8/W2JcqlkMxSjG/f3eKN1pkpja3G7rw0gH5OQh
kMeIn1qiwjbpAH7RJABxvi07AzjEbebGqRyOt6exexV56PQPas9Fu2VfnTy9fxle4pJ1qOfDeisZ
swLu76v1PoqBQRi0nVGigahBJI6KWyT7907kflxEkmLw9lvrDBedeJjZ1vihbnroRC0KjACFRh5t
FDQvHMgpyJKq3V7MV6MW/hk+aOVAAVO9sRV4io8YkX5T/bYeyl4JDTujJ3zk/rlG8R9m63BVwaKv
sm3ZyA1c11ZemQbgt7JmVY01HeG1AJwyx1DZYgl/i12dvZm4750y1aveQHbOFRxy+Zw9X+Cdkbs4
8sZld2Y1Lo/RHRRJuvTjZ1IayZ1HHKb5so1zm7Go9GMsKrUti886zvgyQRouiaTOT7SthOiSk80x
EP4yPN/YjsnL1S/Tgif7JqwQh3L9qM3QafUl5yY0Y6UakEOZYRxCcO2D+H2ilsiiWD9fgPWszy03
gzbO82dSUD/lKfkWdg7GOH4VnazAxLA2yIAf3Ocqqh7+mby7vHQS8qo9NgPW9/bPc6IKb/ejj20w
7NBhybzk/qd9EbHBr4A6DC7azG1qvpCh9YFV4UPukou2Q5AmuVbQjZrwf1t5fK3CG8jY97qNz3eh
vZg6FN9iIwZAE1uZ1Uoho5HQm6mIhZniO3Qnt9Rgtc9iUmRsy9wjD/Zrmo1EiuGsxB2aSbuubrZz
sAfIUFugxF6X7vL+YVSGYffXJ0KuLSotU3YjOGY7GqXT1OC2DpPTjisnZ0klUzNRs0wNI3qRoWwZ
GF+cAWHl027L/aFOjT5z6ZVyxtqPDEgoj0+fuLnjvOxPEsS8yiD3pUYgGPOahuHepV6IKxdgzBpT
CdILk34il4RpJcF7/eJKpzpm0pQlroT9ZldjoPLbNOh0u8ruejKoBdnHqOmBY7CTPvcaTnluxpCk
np2rHypVWXfRU5sD0nTvzCr1rrgSkU+oih6YaYlQRsT8NOmoBEBthVjd8olsajnjxiu4kIeGTFau
TYK/9iXurdKKCTkEDiVSBYBpiS1cMUc6jIODl5atDgLSiQYSgpJLd86+H4dqi3Z9xdNGATnvhJ+e
zbDjr0Q/9tS7YtPpi2ghSQmT6cH/viV2Z47hyqZ4LvdG4Qv507GlU2A+Ko3O+PFvggkywrMLViVb
ZO+bdjervUICl2b1mq8VTP5pLpdLMJA4CyO9os+B2HXI2JyxnuNfRVS1ZeZLRbvdPZyES1wwTIHd
r/fNKW1AadT16xlTX9VqEKySPQCgQNCk7BNM+ISFU+LL6Vt88WJ/MUaM8otztXOOifGojlBGYeUT
YnBEUTVNoEUzq5jGH3GgCfM7hTyL9vsRjOa+yMGKHvr2OerNwjYdUEXXr10QqrX+5v4QB+2H0bZw
9rGGCqDVarHXCf1DHZ3VOJeWVE3n8o/+Q4js6mP78N5sccupketi27ZeVCq24o1UvXPExxZeTyJ+
FzljpMr+vx7E6iZEnxqFHwbUuRJdO50B6rCCGK8UJ7YbZH3MP7mTr8c7wtA6tPmi5qgs1/UHRhvs
RQE3izA1OYf63C4x7vf9wBcltlchEczbVMTdFJQYM2pUt/sZ6z084atCR6Q2sK4bemXKtb0ZKPYa
8idoOLvOJG97di/uNjJv6z7JbVsAtwobqnZGo+xvCs1Ixh/o/dHXE/vQPwxSfnpAlicWtxCX2OIH
CDf0+R+bu+SpIyG0ZsDTo/qfYvQi5DVLMhxXnIQ/uErfiRJNaUA3lvDD1bn9NuqG32BxROgEQNMc
6UcyWp11DF8sRCwb9gSIJfKCdu78Et18+znJWP68iKGk5LGSFCycWO94/abZ9W+vOhCGzK8YMPpk
faMJ/fD4A5MV0pIWRzfd85yLRkOrkhE4vvssPZfVXEyYinn2SzO8OkEUIhhhmYPrV0FSjMDjIQVE
nbaoT4jimIBxtZOE9gPp1U0j1X2azkkXw74r5htpkD8c6BE0QqwSvGQ0d4ivV560+zCrObFMmql2
mkJUz4wPqFDjoIPpvhSw87Srw4t4cvzPPk9lXvtKpfMsAjHzefisyfvYMABnvVH/LCdAiIwE/ESZ
bhxPmbKYFKvVaWoKys9y0OY65hdqKeBTJoJGwGyhbKQAdRDPBIZZ6KDcGZKNJTU32nv3GcKZ7Qvu
2VE2RjUDE9Kr3xXo9RLwmnD6YhwU0WsOEJ49NQDEZTZrqfQSt/C7ygT7p/1quJXGOFT4MAudJ0Jh
nUeVbjDxxmRLfPEpMWTAFTppQ8jp1dH7b3oHP3ZMMoPjr73fcGDuQweVcZuJCngKpyjF6QMnyZLD
5IXaQtHWCYU1YiEfIXfqB6oyEGT6jtk6GdK/iTel2IcTcKVS9Kg0NgIRauGqJnlqtpVuR/p6xODp
1B+8ouWrvglXhu1/vLUZ3tFCp2GYvjuk1e3DHavhQ4wlYL+rGYkHixfsd12fnQBGc0ZpmdQjaxd1
ox7XXNUjj3jnLlja8xxVglhuh5/NU1dlYNWeN6SHhOd0bSwkVuVAe5wFF5B0rQb8df7J2zM6qzlh
zd71uCu2GShFpVrrwdnJtHYO+FcDvqtiaotuyJSf6OOEsAoPHjv0fDqUvq43AyTb4Ij3ZsfYAz8H
mPigtRXpxEqeQRVLyBz+EdXTc9XkYX1zN8E+U+jp04cvvXH/tkY/Mq33ZRN/z5grH8JI/jP55e87
3lvDzRwboCprpPkwrdg92Q0TOHo+VAlWX1uUHea5MH1hk9J/2X23tZ/osVAG27Hsy/9q5jAYAsHQ
G5yD1I0hlC8J9wocf9eVFuNxbrDLwgPm8Q6xHTcQemi62DX0bXgX1vVvVR1wNnMT73NV4aqARlb0
mOTjqeQcdFCwelo7sDXGJ4ioKILaWPKLZGpwHGvChXcFeZ9lNm1RrZo1/FCLNJI+ZgRn1lmnETvG
s2enTUg7xibcSUj81j1WSu/KdmGyiCrVQIRUduBERTd5ET79cSDY4vmLn+SSARA2rItfW/9ifAEk
Zs2y/FhexKoC2psvDNstgOxKI+Aj2WjfcNnpIZ0Rndt7/i1t5AZ628sdRyfGal8YwIaMz/ApeSz9
Q/zLbfCBjgyL1xLOnmgoRC0n8eXgvExV1/8EQoRUPMVJbxWsFUX0qDm6k/CSoPuMtkyABzSAi38+
KoH11yrDgp8HZT9oOfOF0SBwr0YPn+uCyt7tbZniknUsrSm/RYwza5IGLjUHg7Cka4pXVRn0RpXl
lSrwFS3lHWlhilfSg0E1OxWfr/A2bgJUgpWDO7C9VuTuSntimEx48P2nLcNNuoFnuvV690JfsJX9
t2RBLhotP2aQ/4JPZb1b+NB2gjkIzCpIykPVkmB4JB1qWPVNxpcuo0LqW+ufAxsBT38kGcwEl+Yh
v1PP8xkPxOkJH+fV/+94+lV44h4JGs7m8QLMHKMvnm+ZomwSXZsEzYe4MZD2aXOEDrBnI2N6CvkI
jBNLjfJ6jNhVdsUR1woukKJmAY9jTP3c+DgeOl1LnTJ7Huj4CHzlBSdOAUt8eye+ZVM+csntOFQJ
Ir98sFkHr6GDZ/fjiAN9KA063iwenueOxWz4eWFiRgBp2TKiBPplH45Xua4XvDSJ9v7gAiLPL4S7
JsGygDMqQwUMAIePTiQNd6Q3FuAj1k415HSmsFi6pXguSqqYN0hS+SQ62TEyeHJc06dAyWTYLDcj
IyEgkB1umlpRsiJ3QaATSbCYmjsptZiOiAV8MIlElXGjQkDQCwGkg2MrYPIKljQ+V4RKHFFtJgeb
vK/+gnozYGC20PLrPAqVebiY/mjXS52VaSdd5Dae5FgXjmjKctIkgWx4fH/1u0LTYMKlL/cPCCKs
0Xw8mV8havEvofvytzJpwU2hq5ECyEL+47S3Mxuzau/SdZqaG+KDc31aGBZdH3+x5H+dgsw81wYw
Sp85ynDXq15EIu0rQreQiwog0GQh7b9h/KSmzF/2wtVL++Sfl3lhfhD02KgmqE/kIijhP41NnFgn
q6WpK7HsetMohJ7hHs/q1KSTpl8OMHrJl6Qt91fZtF3Bn0ESbZ4t43/jOH7Nt+I8vUXUR4AibH7g
4gCwvXnkhBwY/gNIPPeZEmXUvY3DANGkOrIGYH4piTSdH7vF8Ye8iRru6vuR8Kob972NDUHq7MBr
KI0Cj3ew8BgDj8uOPBtv/HA40XLRtZlJpa+jTMSh6GdC6E/zOam2nP+PDWtBEklJULuVOrO0C3FU
MADMW08JVU3fddzAbGTuX1jHqapTyASJ5rRo8GcbOjCmWaULpNwxJFQAUVPHWEYvufwioxTuQbjg
xrFMgdaAXcNXjT63bar0mbW2GNxFet3jNIJpc7a477cUUZj8Gz6/3TXo2IT7aWSdTnlGEYWqdtZt
TA22mf/zExVIdq4n7F8CXXoDBq2LOuGw41n1eG//F+2UICrUKaEiUTRPe3Vy2kGmBsVqUo3Z9d+a
z/B7qJ598XEmvxoVpuJjdIc7uK6yDfrDXkJ+hQ/J4N9KsF/9J1g5Uf1X2PJ8DTNLYJGhgU7POpSB
MkUW2nC83203eJM6nlLDtAh6ZtzBkLiTzG1oSnKkR5fC7mEXp+MLbueWtyMvBNNdT6DKJIHx/Dgl
GHleOEnCbiwYeD0PN1m1+DR/bLD8Afo6vmUhWLQb6K6uvaSxtf5UBWEByuSUJn+6K67QTgUcO59W
I8da8cQJN2uguvbLvk+CIXx6ji5Cz6kEAaHFIw54ZVGBIlDRDBC+kQJuR/4tDD0bsKY2Fs9Haij6
t4byL8yHnw2CZAwymEZG26OVOsQi6TinWgv3xbE82TUbE3zO7opq4gIsn6TuFVwMiNqny6O00zJ6
Mzp+OK+4kDVN+hH0UKhQPYmsDetgKjC97sYioyrGdvIFAXN+R0JLtT2PxMwogv4Ewd2/VWlH2nU0
X8cvAHe/7R8cx0tA8Un2evD9lyAccKLh1mmyv9zUGM4bRDGNMyDK2JZun3om8pg/QK4mzClmwYvb
TAbcO7KH1ICV8kTo7PKS9EnHcSd+R5BV9lyY8IvJCNXk6i9TkqAELCMrxdFTtsSkKElUeuzNNUQj
vhQeWzYhouyfSLTWA3F11qfJxa5DuxfZxlIt48kVEfXzlWSS83eYCXDlPeAfgvGjoJ+NTfepCAAw
jvUxkOGlwsrEXPILWF47gItfFAfXyKKHvNydvnBdTNMTqxX8sSnNMgPFQaGLma8dwNA8LxY8fSTZ
O+67TmZ4i81+yR6CGbkuh+Bc08IN4aADLV0D2pLjYT6GTqBJGYHXMX+LoVGL84HIZ4m4LG21Ybad
x/2LCKZyWKjHzW9JYlpFJl+HhcdaK/008HF8gDpqoRVAQdg+NTKaLAw0gA3V9k+os8qUUaV9NkMc
9vCOFDPjHRgsze0003Qb7usuu5b6tOVIGqaiQkjtmQkJRdyzIxC7ZK5RLIzPUXZPJXknNPWh3s5n
4Nm5m785v4ClyfretLTK1jFy3FInavOyCnPJEhwdvfquF4+fgx8cHJoOHoKNqdPmBCjI8lI5i8Br
xpjrCBlwJe+OVwmCZJbAqBg46H75p8z2thVXAjGMhmjznt7fRGqJuZ1iop5UwbeOhxVK9aZfCiPC
xRtkOu575ShK+F6b9jpuA5VCyroXV7tvv0GUus0gVEktKe+I02lKA8teHJmOdYImc7gwY4TuQdob
0XoUXXCEFuwYig3kW8WerO9+SIoroxwGWMEkR6ohf79CTs2fRKmXtK4foy1QChog1vFxZhSG4UFS
YM5EH3yNn95SNCBABj8NJoRKNi+hOUpZ8i+cqDBPocXlFb0/McZux/JUeeAxbAzGlM+JcuUtU1gk
5fPzVn9ZUXL01wAfmJiENFaAfjtk8ks485EIsWGXHj3W4YkncTveSrpuSZ7ZjVYi4AhjGUY1F01L
wA1zyJ+EjmJ7L54yeUOM79pofT2XT0mE/XZqaMwgULRjl9C677THKGMjh8yr1ZKhJEJlsuj+AK49
Y7VBR2sesijPl6n6sri7vvR694VuGREO0THqNT2bcJLFyus3TXhVA3mn9y128gSngAuYjqdQF876
nNddSw2DTMpHOzMr9x1IyScLlZtadYo1woWc8y+V0CC2ydDXWPJfJNgjt/s4rsD0L0PPlCWVXwKq
lsbQimt2ZPuY2CSKaeB64tA1CKxyspmoZL4AQrUuP570rer+g9wEMqD1qie2TVS+sSjtPfbDaL4M
TyolwQ5bxJh4jWeKCZIbdZr5APGQpEJ9ucjsLmBuE3CPdgZedr/Z8bGBbuMtm3o4LcoF0w40DbeH
gV5OjHokxbtaTXs/hyb9hcMCBntz8cW+Roc2tSa1krOUc9CD46QwFQ+kKdtnlMR/qGvLsJJG/0eo
CBDLpwyZQv8PCLPHlfzT0W5tP+PEH9CbC15cwBJj5ilcGk1PtaEa4lJ1z6MtIbZKSnWnGwPP1sv3
OEd8gvSm1w/36mrXUCufnbUV4zpBYSsB6z01zpNvJHXnlmxEckUAjqrr/YFm0jbJOrQEOXAyFaq4
/kWFofK9MtTCs5gJby7hRgaNv4Kp7Ys9aGSaI+/x0qIaKVdGbOcXtnnO6ghDDVKjYAnZASwQt/yj
ui5OqHWOev+ENWYSCrdbX4g2f/SgG+21hM9BW6Ovek/8WbO7vvgVXGFdu4zsMi1j1WRJ6DA3MC1n
oI6DCfseCFTi6rUrvDvdQqizYTQ3Aip8IOF1BH5NLbqaGz7TyzVX9TgVy9OJ1a4f2sokHAFc9K5H
m+36u6VrPe8iKkBRAVW3O0CLrTqtMardZvorVvHlrdFCPKJnp122KXy1+wwutzjSp95tAyHJpSQI
KmFDSob5op2g5oIF2dBxkDdn+Qugu3W28ztlTDwLDYbm/rA7I49jWK73WAHbpsqjXCQz3sGDRese
9Eca8GM9xABNHH+e8+Y7qxEze7mbX4Sc6JH3V68hBBLJNgWLeIakK6eJPGvLc6nPLIzvIUnGX49x
vDbttp6DSSyCc+Pk4zb/PPOwWRzxc2Jej4FFdDlCq2jXH/UNvj+23VxWGljHzqkaKHVGuWxRkLQh
IdCV1HkjKjwLMKmRJBNa6ZrSNdkMmykvOuFCe15Ih8YX07a5Bj5Lx+wVm1B8yG5Qll5biGYdwACI
CifA0vJ7hyCgoWEWsf2XZDTHiVvF4vFHbmDJ+n54S32tcXp5OqtHGza9PI1v5YMrQGgqCD8XnUlO
t5DCSi+V0Z7l9DyOHB95Xa7mUiZGpDoXC9w09F79vEEAavvVaIhN/vRTM7j3JiiW43Zvnwu1KU9S
5JxO107SYuWF+blJ8A8vdOr4oHO0cNmmMct4396W8iVkVbqs0TGMZkT0kxX+/Or99zAmSY8qlY3y
icG/RfjEl3EdMN1WyziZukWgQYCW1cbLcpX3M483dJ3f+vaAYNbGesXe4N7Qtdfi7RbQeARZWULB
mV7Pfg/1IqXPVwEy1QSqGea+r5xvDAofdAwUVhUcgCZhlOUkCTxKXdtCv2AMioKapVf672bh35Pk
vBiApddA0Ycx++NqJ+T0c/cuLYrHq9hPhkdzp0EIhDzKbmfIxYZGGtsEJLQihaRxwXzz1KRxWjcP
CPK83SCKsEmDdwKE4iEOfVOyrq2p9uk6nPPv77SDLepiBz3Jv1M4XzxRyjK7Hjm1aDANi69j/DkX
YO7H6e8Vue9/tUaFJX8RYtj1GBmu2SAOoFuAUx6RbiTo2SVMcwLEHmUU7xT+Swdykj+7xUdi+H50
1fLFjpStZSqeoHOz9+cCmRV52bLZMKcF5VVj5BubAO1RgldGUYqJ6zteS4K5rI1uK+/txJl+gHRi
HBsKtS0Z4GC2VZQ3r95coinRkFlQedsJsh3tHWca/7SY5vsN9qlHE8JA00dnVibMq6JznwviVrnz
jY4+Uw/C8ufGIZm/Xb1GKEeBmEQMhSoHJbzW1TnjXYyWNj2F7uoAzrhtQFgyD4IejQ9qfaiLnixi
izASgQ5kK4x0tLKpgJeTGsnpKsk19GwNMB6IESQhFvURR4MphWXrhfMuhP3Y8hhvwbdgK41Mulny
yELQuvYK72GWum1saD5Ive5eX2BRCM3PWMQ/lJM8v3PRk28aGTg/AzthEbzoom114vhq1xWiuXAi
bsAqo2ku6NNl3bmWu2iq+UhoKTve+ay8oB4y+o/Etuak5dTNaPE60KV05u3DiCAtKDVTyA6Bz68B
HmZIQSHi6DxHwprivxdQd5LraxRqme5wWw+RTUfPE80TjE9Zkgh+v5LAHT3j4Mf/mJ3crdK4CcoS
+oXOETYxWtM1hgsMRXxlxwyCbcYLA8GFpHJJP0Mk8nPbEDKvQRJiiG43KcEzIDxPy/33dsqCuM/B
V49hgSDOS/7W+Gn852ihFWDNXnmnrcgVC2WTylIxW0UMboioaMw4LEtDOaLrqegWowOK0soIq4mb
4aQeV8CE5uzvQqRZNKgt3cX6KLEJ4DHycOhCEK8J5G0+MVuRmxEUDMYdu+gTDpYHePcco+R89DgJ
mPPSBeXqO85wIvZyeDefUduHmK5j/ExqOn1tDPs2TeNh7GFKzkumw+xKJgo3loyFRaBbyEtGyvAQ
CjuVPFYYmsCKmnXbdNgQEM27Gp58VCI1o4KoJsYED36tQqfqppAaF3jCIgh0MIu8NBujDLXSHcrt
bLDrzBqpXlNub8OqHfNHVbbIvu1U6mIjzFR3QBSMH3nN/KMnFy67+l3EepxQa1vnuZ1OgCdzP5x6
zU6DygHukSRa9btlQO+5KPDYe5i3OLbYEQeD45+zWHRPvmR8F7RZSboWsH+yDViLk/rLE/GhiDav
N2Gl5/64Aslm6fsHXy8MeB97YK990uf6FACSCvPikMqawUGAuEA+eiC7S1GYVyuxZwFuBRr3z4/F
sDLT6mGEx4REoaS8f+Xtw89TmdsV7P9HpOkMEN9WjEL4LtjG8AkjEuFG9/VDDlEW1Sj/cIkdlkAv
vfwek04q5kAp9IjH+PboI2IKUFMsOiBRTFz6x5VIRmyw+2ZfYPA+hH+SGHWsTKuoXn4OrwB68wPf
7IFSvCk9yNENE1uW/nlHpVBHHqQ1M7CXOiuuVV9L9B7AfhJfed/MyXYziNvnpVrxDL0gENuDSmly
DsVLAnNphw5UJwjVXoMbC296GR9neFLkXCyJIR8nQfDtOCQ8WVaksIL7NBfj+rfF/L3cRYfwxc0w
A54qTnxnhfODxtAH1UCI00qUyDt1FXwBcHl6EUf19/JlIIdGnonyLWcxkyQJOuCFidQUn64t0dBp
6U+rawwoBxeroy2IY6RxGk8s7CcHy8tUiDvJ5GvMsp+BOYkPsL8+qFQfLZ6Im3X7zAdWdQS/uplc
I4807dJmeCJXiqjRfSQIdwFrgCZw6z00AnZ7kZr99DiuasbW1X6D4kvq82dLTFE1ylp9LKHxGl+U
5u4cHRBfS4UaePtCfpaOwf32ACIhKDYjQVMjADPdb4wUjr3/n3xbGlHNGYjn0rStRjZO6aNBZx6a
7RPIcRTJA5ymPJd/jGLHptFFG6JzU/KbkOtN2ypg8dVgz9TOYQjLRPRRuaI2GoMogtW3gwdQy4XU
HizqeFYBFUW1W4gY+1eNTKFD9UxQO4gc2JPNb+UE5ML5mA0L/nsVojBf6+7Z83Mc4SFYz0PGZq0p
3KC5Y1AcENtn20LamKDX+GYaeaMKJNUh7Cc+ytOGsDZJuUpBkkTh0eILsqrTiBzdNeDwzH4cxa34
akRCrwWvEbWqctuksuI0u20nUzVpf+2T4RCcv8l/hd8GKYzA28R4UPau/uDAz1OX10O9KH9zXqh3
QUqm9n9ZadunMqLdvCEzMmsQv+T+Jgf94fpThjI6Qb38wYd/7niQNSn3zCSUz8h41p4ZxHAeSyH6
rw3Bh1FABAWtWctiHPniVD7NEwJuXSzLFHnQCnZxv2IhJz/MfuJcKBA79t2hh6ZnghwmjP+iHMIy
TtzRBK38BW+lWwTXPq4Z0Rs1PGUH/guYTtFb78I8kCTPDn4SM+rVupVGvdBPeaAWoEtVLg4PAG+S
cJHipv5J17pBls7OenS39yNXipJUQ6K3MMPNEYOX9F0tn1g6w9fwxXQ9SKN2bY7Yn87+lWEk3/ik
WdpCgjQ3DnW0omN1+G8CmZjYBn846kzj3kUERrv30CepDl9h9Dvw2nQH8Wmlao0NaKJbwm/UZK25
Pqlyt/QAim2/yZlq3/cP/K3KqfC2DE4BGB+1cBchJBLEocCNiBPj4IcDpwpp8s+KtStaGh2P1UFB
JmKitQ8UfSN7I2jRbXv7ex5X1tOEFWJi3RhuKtf9wPd9sjRC0vm6dFG6tOyVB3LbrsTGZ2CDJjUm
HuvyzwHt3adfTNvAWMp3nUeNN2CgbG+FaifmxniR4LVaRbbfmWzL/a9u6+B76o68x7Bbbxx1QByv
eK5GJ9HLT9q9/tMqUCh6mk8MG67GffjisXWPvk7NIlVrDk/9KYsdbQf8Cs8qEuwNyqTgANHsxc6S
dknHzAn6a9iGEjaUpEmHKx5tzUaUipx35EUE3x2t4kHMnGXiujI5dna4ZbIBwdf2OWB77tkjxpvp
NxZIJyRewmChE94dB99jVJVLxN+bhV4KjQ8fnk4HYEKQ4pmgMAfy1lyFoQOvWqEjijfyefIFP8tN
MHBC8B3qHdimMpp2iosTNhwZbZo2I6JFN2a29RpaCVrTmD6HFj8rvHvdySEEsGxktoGL0QTn96my
QFdPSLFvNet+UvCCDvMtStkdq6Mub3v+BzyK1vDYhI4OT+ocskPhToAqldpDAJATJhJADdjBV9AV
uDDLQBJMPf/i2TKyJgPskmAQLF0f/Y7MD0iv/YhBJkwYX/t4MdmjxaxuBJdu+kJXRhUFkMGhkohw
LxZonl8ypOCQZ8CxWxGPzlQknjqM2PxKj9Hx6ZhF4eOyB5Xm6e2jg9LYpD6fEgaOFTO3pa+dpBNO
OfY6Wh4juTAo2z19UOz1TNVs4H0XXDX6+A00W8fQUZCTt3UO/SZ6m+f1D/ydufKRhZbO8yqbsrP9
xmYOLhAaQpDokX3myDbFyUiuvjIkRLgDzTM5Pu9/wUqFEOzfHh6rrJGoC7Os4E9OI12nDA9DlGMw
lpzn0Em8ZboVh837SzrJDicsFfdSj79sG5V/au116AhadjlPzd1UbSKzHEt5Q7wNbrx8kRitUPsv
lKi5+oX32U0RaBICHNppMJ//tEut3yf6I5FiDJc+ng+OeXNVnwgh9mzhujuM9YP0BI/IXuR6ANqL
+lLig+HBsy/ns+kTzQUTYWnGJwV8pgnXqEfBuxDswTV0tpTYcFIHQb2T++NnJHVwsMRcS8WVb9ac
oN7m6segulDstKQrBMOBRb+V7YFQOfcnS6kW+86ZfQLwErldwdNB8PPgmiMGG5URyTYXHaKjEClN
udeEexnc7M0DjtekOZZRuAeIkb+e0K9kEBUwPjtxfXGfYwQC4YGykYXkZEm12wj4k3MlDVcG74NW
i1wzycuVmj6mfuWVQ1WN3purz+FYRzFM5M4+IpsTmeP1If2i61Dqnuv6jh2NYVpYjNIXCk2BWN6h
97EPMj9B26iMSVG8KOMRoUIRSGRm2uD9xeUhjwumZVu35MFHE0nW4Xifikq/ITF33p0rvMhungWX
l8/Qbz7l5nyu/YYUGrLjBZLbW8CimGr0+YL+2GfrEfy/bAbwK2eIg3JKyRurRzHqmmIkzSYDsCZc
IcK/2/3njzP/H5KJthyKrTD5wLAw+p++jcK1HFlHP0jECUyh+ShR1LseqlPtPVUqNdbpspLuXI5A
W/T9nAjoQMbB0R6sIC+UMkzsKOBKQXodUAfcNd7uOIyeejUiWMqM3g80flYM5qFEiovJmH0dmadh
ZuYSndB3+8GBDonVFDJ8JYrymAzdRx27NvNwJUcQIWxkc60TAx1G8vt0ZGJg5AgteIwA6e1ReK1b
ns+yu1R0JmoGQ2d/x8fy9806xzSbaXqAAbKDNcFywPPBTF5JAXI8JC5UjqQxv6nUBGQsCrJVWUs9
2phWAuIDT/gyRgtYDQhYedu21orZShyS2HGV0WAMw2O5gcVgwEPSBV9XYR0o9akyxA+kTQ7Y6JW+
H++0q7YeUnKYOvuwtymZWePrIy4fkgjmXsAQcRL0oAnmSm+HsUjHG1ud6AlfgIgsuRDfDrRHDylb
4qIl747tUVGU39cPpRA6VvsXrg8NEGOqyA5S6jewXIClk+HuudhZZP66Q6ffb2m/PRunjZD+7Lof
md92bXc+ylvsxBjNN/Uc8CxC3ZkjHmOailVjTVwECdMc7fkJzyAzuU6quALC8/5LRv+UZlw4HsUt
GzfW7Ywkligju6VLUZQRImw8Mvmj6+tRjE4PkvUSR88dEpZY/xebhsccS19X+OPFBgADDdfGmuDt
owag2c0VLlb08XZfiXdD9sYv30qUQhEbxyQi4wYKBA4sBL6rik3Cb5STLuHGsGbzy+QNcIdRgzOe
X7aZ1e1ina+3dtwMc9mBgNXDgVQ/wgBS9fRVw4YQeVhbv80ZLUd2TjKdE9KW4jsZp5YggFIvz2QX
pGXUDT2442cB85i9K9BLzfThuJzZtEGPGCFY6B1P7gh2dEs4T2ZWUn5zEGG4QXQbHymW8+LsBnnE
EES9uW/JKGBSS1P2vfmejKcv+oxBaGpLUheFRgD9Oh+EIRJ9uMgvmWOdrP/tX/eZJ5ZMXWx38mRD
T+PnVLsRPahYKOjWL3cCqu/qYMnfMgHB7n2K4JlRGCOo0c0u8LLyvp6AF1+W0tp61oxuotUoQJqM
mzzfEN/eqaqxrobtzwCBies9XnGZeJ+IqYNWYRE9Zfuvub8N+h+gFzqGballw1F0Dvc+cAVt0gzB
EScW77CsNZl6OyGIHVbHw06uw2FtC6R3Wg4ODmRLmVUHj89Y655+4Bz2syy6lmP4YsEJs+F1G1S4
N9SsgyrwvM5AwxqTOPot2FojZEj0ZgAYLnxAvMkfKXea2glk+2SH/7K366iKzhrsKGh8tdin6hAG
uW0rJbLcS2HXZN3l2qfJHcnMynL2s037NcJZPKMz0assRTdMaZtLrzfueRDFAqmOEFWGpYCb1RPY
e9jfsa4hiUvR+1GfIdobEZQVrqWs55Ea9nkGyiOpqNHxTLuzBFIGGAkeFolii3X0EKY5KAqSNU0c
Fg5gIfbFTB1/NBPRZD6HwqdQGiSR+2TnPRyMcNqA57ANZX7gAw6E2QhdYQf4iA4aO0W6+FWYoDOU
fT/HYe09amNgR5Pmgsr/IrZj0hWEjAs3t60qC4AyDz6aHAJiiHzcUTac9MCq+Z2GglAU5zGUSrSk
yCJxZ5ugYDu2RcwrjfxBWTsNJcSzjp9JJx5lk+FFMQdEQSqjgK3r+uL43oqGN4r2Kat78jmPZL2w
I/ZQJ7Y8Y2FPxnuLN5giTimfH9gv3PiiOizky1ktcqypI66MOWphDOMahaJgbHArdso9uTwcKJpF
IM/0CGT1hwsmatVx+MOU/GoFjCRxe1qnrJGch3i+VUhD+O/MRWqeWi47TUHk5QkYs+2b7F1LpzbC
o+ILkes7d62RthJzlMUpRyvRbq3OEK1lx1PTYn/PyJdpHkPFI8/LHAcvhExs7MdVyaP2bw5/z+RA
S7rjVyYngUsgn4Ia1A7tDltUiM5I6DMhKa9fs+vSpkEneerCSOYo/ho4JU3GvAcQvGtFGJsTXsDr
QPCaiSSwZDw+IckafGJsKC+ae9MYbU68ch1pnKJIglwU21VCt89fuB0fFsdu2AnnPUhlWIY9pRVE
oQCEHy0YaPXw41zSPvSh7PkaDo3NWAzIMoyHIacuJ0GIb4V9AakLUeqxqegwW3765VIgIwvZAoRd
NwaUOFcB+i4gOOxbybvt42kRu+pD2WX/OvIW3xLMV9p1vUe3GAlzmZCbc3OA78tIv9aXov37WXpI
vGlzjJ9kfeT8aWuT/E0EavuB7eTfYzedJoD+meMCQx0gB77WPMbPRjf42S4l55gXTKXePCpKZFhE
B46zzRAUlYVRaGkpPDlMiVcj6GC04VF9H49Q6OnULEshN+qWV+fYq3eREkCvOrRqK21e5TTfhFu3
v2/Xor5vogwsqKHu1rEjNXQvkpPStcYH0ScmbRXKvguWCrcc6S7dESqrYtTHdxPiTMXWc/q1BVQQ
6CWAKGlmFslt62QwMTjewkI6hF8JqH6f9ibsvjyOFLKr4a97XQ/jIGCSRabcYLR0dok5RUAKPvp5
lGuS35m51Os86ArI/VhYNGLsQWSUA1VJ0M9slHp/VS1vpXckIZbZEXSj1YWa+NMSE8Vn1wxPiqxY
0XtHyXkywsTOC3llwiF5wlVa/CVR0jCStRNeUcJJYDeHokNGmWSlYUuNkeCEJMCVoqjReQHrhRKt
Ye32Kr5KIAtggYm88ymXRrTMd8UCU+Uf8ZGYSSjhsht96H/oDwyg/mV7Yyb0ivynnyA6BpbgRMkJ
uDbS8YHNp9OLFr80cCvVVc4xyVxXHA1lO+zYiynLf8SOFtZJjSEXiZB63G+pN79dAd3ipgWCzN0J
si9bo/xPHZVSmG+w/ubLm8I6O6xhGIsrkvcYJp92vj3kq0VBvRW1+ZJCLTKiFURjx3eCuOOzS+de
vE4S4HWgXQNmqyATr4pvMU3qY8k6rPeBhT0fOzciN3uhRNwjKj3Z2gZj5//G7H9FYxkRArfNs8eL
gu0C2+Bk22NIJwjU4uolofJAIq3MAM5KZcnvwhnF9aEVUYczO2igVoDmGBCt18fPHWTi64/pOJAi
UNMNZDdz16WpfPZq+iNXUOSftD9sFJUfAgiLeakFQ+VGeN7y5Y3ZcA19Qr8x+yc5jP0y8CqeqnYh
rohfbkVIVwFBMFPkVRB6NCOSDZ5gwjOV74pIvTOd30bj9GG+oSMrGRaFPEem2567XlJPqwkaMo5y
bLRv+Oh78uLMkKaTqTxxt2G2zZglvEZEBrkwa1SyWy2I3yOcuYo4kUpf3sOyr3AD6VGNddOnNva+
2e8KRqMsdjqQ73m9FZMPiF74F/lDL5T1F14e1eQgnFrhmSdBRI8/x9ztl7e6rcBzThJDcaawLqZ2
bCa3ano8g4ykwqd6jIFW0pksX7uJrhzVPQ3YtfBgjUIpfs3d+yP5hECci7ZB24nn5VRea0cqeLGj
O/jYT3nO8RumvXXqibFv53PTjUE6bSyogEUrdS4+JmNfCDLjx+WrSAJyjExifgN291PvStlnzAQT
QvGU+M6MdulSkiDLwjVW3Bs34epDPZoQ+mt5Eck7cmz8CzGtB6kepKR+1A0YRcDnVHW/DKdslNyg
alsupHYap/uOMjergKINBP/hKaG8a+vZUrlARso6jeYASp+9Y82QjjzbZ4U73klJXHmOmGW51hJU
Mv/EKgiTB6X+Fjk9IbhAIltUQM5x/coT9V70DrdKvqu95MriRWNjYj+AxUVj+PcjSMqQTly919AH
IP1Ii7LqM+hQtkz9tyrsbzwWbDNtDiIUlm5DhWIgug7X9miJyE/+2/t5Zh7tgL/8t/t1uNVjI92B
uPGJJni2nJ1f5aMOK+JbDvP7OuvGRRg+wdr3Kke/sdOJlf9lGIq9zyzWTdGEMDM9euXyvKkU8oNZ
nr+1RU/3vLUtjns1KNQCpgX6NgA0F62bLFYHbWyfxGEOSENv952ZS1EMtoL0iO/QMHP6yRQNHMl1
A9GvPSs+rexuiTejSJ2XQNebWDcrROaHDPj129qLoOKRIu2mynJrSj4ZMCn8TPu1QUVGYTYUcH48
4M5hREBWInjsidivdr3JODleLs5Ag2WaBNYc9UWiAv0hfLFJzhxqfJBZj49QrWz8F9WWArOF+ZXA
bnjvyhSWtNoaOvwCKsks0d5ix3tKAO2jyLu089R3fK5epbi80IaJvqVrkV6kX0duGaamSQrPzCkF
14oWV9QtuEqg0qUl0BbD34PW+swpSAYY7yCR6uKKMz2PTCnOjaji+BsVDS+LIrDCBDZGPazl51pp
/h25bCTuUGhsh0paAV3CsKN2E1l1fvARhJeYvCqsbBEuixIW2e933woUoCCeYD8A+z5XeMgN5P8b
7wsRxnsM+NY3U6auVlZJDE3EiaQU5eDIUAZo7QLbznJx4yQ0CEVDbvt2abEShmmMoDce90S9EmPI
ZfoHVxhOhxlRZt6G0cHsrcx+A12eKMrrMc232eib9Cx9NRUqCy3qed1drLrAOS9i66YVIN60ioho
qz+UlTwmSAbEtZcgS74yJv6MKK0PMN7IfJ4mH9Q+iaaOCMeDiHM5ByeM0yo6c4HJJJvHg8OHO+y7
g/5rZJuyB80+DQkpaHQABrYSBg7ICyC+NjOttNUSR9LfbwBSiNUYkx2E26hffyQry0Qvdt7Nv3cT
hFdAbQfz0Za7ac2CJpj+42M1mGFd9x/vB55zX+IXTYy+/Hd/LLtohFTajjZ0crhkMc44gc1Mscol
cHQfQVxzm/2TtGZSjlHSh/id14eVTCAzjmqs25b/cB9sbO45wvsjoFmxh2Zm4wUmE9wjReNr1uw5
civP4kRbRKPiphT55tXpRpff7RNGyuJF108VAS3F+Q7pwCx6sLu1Oi1TyomDgZwyLbsVUx6ou28b
0YU0AdeO0/iq0YB5iDTFurFToJzsUcSa+8yjXsp6G/VNW/Nb0oya/DEp51e1266LB9pk3hcnp6np
GDl5jFQ5wrhgtZMygC6WZx6AqsO018v1mWjpPBZNDbB9kGUGh7KQpU2sYWN//IGJWJxnwPYP4Gwp
A+xmkNyJ+AyyKH4/1XzI3PAgCojgB8FtFKzDB3gvXY1L7keNjsjZO68UndbuYw6L41gn1UQEN8Oh
sNjtWn+DfWTtNGt3NimWqI55DTeZ5soB5nx39w7/UW4a4+c0OHdEajrjhC7E8kd48IzVfyXmXmoZ
gGsAFT6uuAujHaPoswCurzX/IBHy8pABwZ69jNzu4kU/CfKEGvUJYre6XjvL/OEzBxxBpzSn/87D
cclt7982JGmD7gEaqvg4SErUB3/PweIwjUnFHj1fSZjTJKQO/6DRx9XZHRx6mzQqTkcVwTBS2Uw0
Ouq71WLSyz2wCEyNW/vrT0FhAbWjgwNIXiR7pS72quGxN+aptgugtxoydfCbxdx844FEzr4TH6lo
8Bnar++AW3aPYsFVDfn90oGL1guec6VyXnHZdILeBpfP2/+0UT1ht+LT6exAQBfV6VoU1uI70FVU
0/kGUQK7U0bAm8VG3aTf46zXfRC2osLYzN2CydFOQO3//Wlv/y1QQDMGSa2GaQQZ8MQ9omqCFlH8
Tm0zjYTgqeXF9P9t6pELcyV6M7wjrroD9eQ8KyDqCxVZu2Y4m15lsjtSeK97pylx334DqZNNybEB
eyBH206/CWeUtpRvaQSm87QAqzhuCNXaND8tAyTQCXOavl8QbviNBvS+3E/ixrGJuYP5oVrEgHx3
XQlnv4K8jOEwYJJ6A/+1oW6JRe8hhwZh4VExRMNFiolHepshW0pMqm9rTuc724Ah/HGtl/4YFfQ5
c+OIklQqkEXFIsX/u8savOdrqdG19xpbI6T4aPee9kPhdhvpDItF49f25OiQp29dowoGycP/vEJT
vi3mHYqsDHkh/wKMvmJGIYo9LAOHzXQI3xOjrAKsEmuJz/b0ZYz+XPNrV4KAGbgDOB3WlG7uTi+c
2YUza1o5nq/mUdCBHCoh8kbvvdZVWAgHE89L0+eklklTiWt7LLZJzieUsDawJV2UuwVLyGd934aj
Ek2oov8NWXUbVejwhG850+aoGl83PbHcQ+vOQoqq7vEfuDDFBQUf/4FrtY7nom5xScgpkL64XbQE
wEmmd7dFiia7LqL5TGsvuiRcrT976fthbThQvrUzAmorBf7WA2efbHIoYbBjy4mO44gFptZtZNx7
bVMf3ovpojtMdL5Lub8Ew0iDlm1RHvxYEeizlxl1MNP83GczHeBKp7lj1kOQa3d/8PDWUIX01d07
tkFw8Muu/5C6i6JKlxxKlzfHuGlzgG/Ofoa1FXJ3th69NA3CSrvOf1ky4i8v8TvUFL2NSg9+jh7r
drAgmb12YXEnGNrLeD12bkvfeiLwQoZAXlG855lqXKgRGSBKcLHwR4aaeKfrv6egR98lyUGtGDQl
kbwM7UHZgU1Vhj8c6YnTowcypKSfXUIL63nqTaa7F0lRwByqqowUZhgN9LGDgutvfMnTW9YS2Z3a
m7Av6Y1muBirwwCiltraYsHO9vHGeW4o0fk6h6T0BaARTz+VdgQKTAlqRiHHjuOU6YB2TxZunexW
rK2Yv9FyEvQ9t+KyHOMsK/MXrhZZsNsRL4GtQGZByr3eqlwYlrpc0Hk0T5kih/pZ8pbaFpA+z8AG
VGZ1BY1y89yTm+K9z+XkLDk1OgEDvuQqu8c4pYoX7M/OOH3NJtx6hbSNRA4OFn+CHG1HB/6Xi8h3
tK18i2WfBt/nYNvgoM9lyiYlQjTpfkWFzCDZs963aAfUtotYUwcEHWk632gB5SA14/rRWkr3V6as
SsSlVCdROUmA2VbaVlv52o4mWavHq25qXLKLW7g7U3UKECJRwKpdkfqV6djDLpRkOze75TPrhuNG
gC7h4rTS5ZXkOZKVVFU3qht1jnmT3Zac0BDJDD1T5pJs0SaYhSP577ZLBuDVaPZ/ZNAv1Vr/eCHs
0FisCbX0FEwmjQ1N95La+w9Bqb7B17pTTyxtdG1iOnPWJsZcRsymMmoRyLbCnO8QzdnOK+ksnaeO
Kq0MG01UV6EoQbgH5cOuPhILOxL3J0Kfg56TDMTvt36LOCZ9LT79io0ItpbORzY9wLhtXFbomiOj
mV5CDvDEgFYhSsUXvKSUt/knCvfATT1Qan5EAZZQQNJoJ5wokC867rxdQrhvBo+uhURBrE6UI9ks
yEl82Eq+NPOuGXO9BdZwNn2/AMYV025auvL1DuIk8c3JNOx5chYOYiCeMdwFPRW8oS6lmou3vXau
KRqx6sbONTjSzhKbg1wdzE4wcw7a8qlhXidqeBTsbm48N5ZETeQs+tygmqu5G9boDbSx0O+akhGe
PL99rdH9H0mDSJXgPejJjtZI8smrG9i6v0wV6psWyvMZiPM1V9kbB4eb50I7aKhs29yWAj4+BoeW
eUKBin1e2PYzbHUuru6R6FnfrBBvggJ216Mr2NbcTjk3SIQxxxDePNIWZMzJczrn0xSomVaDgmFp
XepumnHvaA31TuNjKnjHwXIw3Yyjyixd6/XMtntNEhCCYC40uuAErBP6/8xRZLkbhLtRdT85EtBf
rkhHxeflh/Q182t3xfEmqPA9hilO2P1eaGPDMROoJcSlbBEdS+4FrzJTzZNkVywl9QMJLn3jDLLk
P+rdVQnK5aekIOwm4KzuAmOxBWqPunv2HiAwdxfYebayzR+XT+uG31zVWCr2zPBHN0kEFxTY3NIE
4K/CHhV/kyZX5YwLsaDNmA1Ob5GotAcJveCQho5/RBQHuMviQNIlpPKx0ZX/OeKV9hDFF9PY8reJ
tRzvKZec8CGWf0ohttxo5kWIYKlM6WkEXyRZiYXS7NnqSTXLz8L20SuOXz68wi9rpXN35zN6+ym5
tGgpVSnIkezSqhgGLcZV6I3mYyVEFPuaDJGnB1XfZI/adfl8hb38T2TFPX0O6sqcV6khiL+Hz/OQ
bBZMe4WXPO2cUQt8i8PCMmckQuvZQP8Kt1vwNmssbHmdg9d0lSRsOsLFnfOGXic2SaMIS6VOUCrR
uxKScDYWDYoYBXzotnR0tU1BmCpbIf7IUX1eyITiS5MZpuimWzy/GxeasYPXzeHne5J1W3imboMm
Uf0z9/pDeY2Am9DG0c4XA8TaKFXVRJxaEVdUSd/4A9DRmBwINNsSq+7IYBVJe9NNMzxBazvY4oCB
+v3Sk1vUHb4Qpy2P+7h7AFREuJX5i4ky29oZS6KwIfAS91QGVU+eMLqvWFvORJryi1M+KtAzynar
OdpwlTAX7Hg2IHr6HIK8PfV8GpZR8EmUjlJcwqJ3h0nzCvCk18VTXq4QIP8Gw4DVO6Odf8dPwtHo
z5iPDByZyAFN162FKWpjFL5nDMA0koBRwgjDP/v7IWskeGM8VTEJIgmrqGxGUare5XASNC+nfS7D
pkFZLP0FtzsJZf1XkNpqRZsiRg7P4O3UO8bEBw141fl0fdQ33C3ubije8q00q+rc1PEx366rpO+s
0wIHfzyzesStxbtb8qma4bkdIAd5iEYDz1tLOT25qFASamrPb/G0bh8U7YriBr059+xwUQKLlSMs
Jwa5g/Zb3QCZWRbRYVYzZPpLwsITkVJjUXoLb4H1nstqS7amYjwkDgEfA6uhvaSC3yxWjAQSLSf1
hYVuVCEqxORnOj997QU4xQC9z3ptl5r/ALL5nOxl7oqdsjWYP7NQEv39C+HwLnnagpGrvfjmnSML
Bq2nBfIlt85Hx0DpvH0HiokVLitbiDKYEJXM1rKSokizSS5NNrGri9PMtWmssUf66CoKzAfhDJ1f
T9ysAf1ReVtytw9opzMUS+WtZJSP4n2wAwik/dKYt/3s0z1dQcYBkjKPw3hDoGjvES7smYJBddDO
seJWa6HJn943Z8IRKcc2mnapzePTLaYpRn4/x45H8hD5lDRtSXnhU7sWrqYxxS0jJoCdLk77Gbey
jviP6nDYx+S9DzzL4VfpSRh1VECR5waLwCYulorcyLE4JPcmaVF/lh5j1upDJCfAoN3v1nK45opK
F5zB/vYkhG/8Q6Xtifd3w+PtZ+NyT331ILRkBwZCqwe4l2tVFy7jAxn4qnIVlPqV+QOcyCGBob7E
cG4VoCtLa5N7GRuRFVySckXVHLQiSenkMdOkWVMl0uL0oVfmU/Co4dNbXxOBFQhck99lq+152Wcs
0HKzzzgbs7QP0PbpyuWPMV8usXdNqr8XVQUPX95qZCfzcEZT7tvILekO+ubV3n2C5488X+Lmh0Hq
jWTSTkqOSom4wKZZfpCwCgpd11kWgFDLDsBpN+7QBjPQ6LsYSecL2CBCDpom0/JtdTxnWCxpp+zu
uTRFtLNjOFy1EKPbJS3TKRNetTMUc5iXUCD4/C1itNrxCsVRv6yp890DbC/qaraex+IUDwu1fGS+
aMUUIsJg7rDADi+xg9QPKl0y7EP/TeOkuHvrZG2p8GgdlgT7IRMBfs8+OifEOPKf8azSDD5oPAoE
wN1XiXfEh2JKXoYVh38cfBe6pq/9eP3KxIGLLDPP4AEg3UaaSpCsnEpj1P6zovI9IKKFKP5VVYMY
ky0p2Th/klAnh+aHG/UvKI0XoGM0m3fBMvqO1ksNsCuE4sr/lJq3RFQyuAfM99v8dBdyGDqpUWl+
6j1LRaW12LwTgAADpmTiZaAP02hj4kSrEFtii9YSjfD5BZzem8xiAQoZnPF1009pkxC/hfBE5ar0
x+x9nPsXKW0KJ9oQeUPkfQxhK7cMiR14owGuehX7ennzYn+J7a/C/OCa/VkFdSyUdvwquyAcwdng
shl+znKI9QW7akA0HfuvfecvMA5WlX/Xja9KPUPvWQD3s687A+smiR34bAlGDyJCwxXf1NYqG6Tt
DoWNyqEcW86QIumhBgEZxcfseS7feZPeS8J1ns8lLSwcq2ATKNRnXCzqPxprcoJqZOrf/XisX/fY
Aa30xM/eHTm5jU8WPDPLScWGhXG55lQ1AqGJN5KINQIx9/8/DD5m3uDQOmAWK3m85pCABsu87vVc
zUm3lwuu3lsmmknqdfgjPEvvM9WDIlLP74RJFQ3MZC/Hsl65uEXKwP8ong0yVLlMIhuhw2bwkcIi
Xq8KFKH9dXBiHhzydHVNsL9JM6EKmGtKp+fQVPhskU9QL5T/j/Pwe+cK4wd/CW47OTEeSzGW+V8i
DOlgtZgkpIyiUVWCDQfhA+zORWLzO647q5rNyfTS0AUAZaPJYshiK+0Ve3DwtMBO0/eC3bX8sP5x
xjnr51NoFVbTKwCZrJ1YQsJMgtLzghxfbkPEoo8w7GKpViUNYNnYx/XW0zQKY6HG/o7wuSc+N4t0
TxsduuQCR0r9SC1Wm6fbHbg0UZ2DR+3Dp9rOKoU5wrx1ni9TM3I4YvANY/rLkHTYgMeqReqVVXlI
Temwz0xqR4358ERuLejPXcC0Mxzobl1lTLLfbQjRN6KYzusBnkkXc1ro7UKUiJjvs2LHl9OO0uHc
Kw5fCck812m+Ew6GRBXjY7mZFXWsQiZxMi9esdo9O3HIugDcTE3imHc4fmCLubectnZXw/jqI0d3
kGuvZlR42tqQpw6WB0sXnIUG3ulSj1v+wFFUm/B8u84GlU7SvIP5e0TKDGInzf3lda3IEkNzuVcH
X7+FoM92/mp+nRNLjRCDg1nljo6Ks53Cz4wmU4dPr3vxq+gWHotqWn6n23Acsyep4BC3vuAHaQyU
8ig81Ru1g0kUM13NennAoOGBZK7pwJl7DOsLsI5FKs+SuJtRRCyefk5m3dLIEpVe2lkrHZA0N7YV
PCcj35czK65PELxgFZiNren/KXsjgsBNB43F4/DFimLnsnizhoxahFLJA4gdkrBMAdAahV5OOS8A
0O/s0Q2scWJ2uR+jbzVNMGdJxxmtTtKSaWHQmgUBIptvwadtYRijotKbDrNftxLJIBmbXRPhuRb4
mxFVGJR+QMH6q6pSr3StHydcYycKUAFhIT3E+qyZhr/clTXs3NBMQ36uUcMNtHYipkhv/YJseyik
eBomwZA/hUUZmqLll8uvfX5eX1sRb8g5Nuh1cYdqyKz9EB+UuzzAZDouKLf8O3EZ6vR6+CA4cv9g
iqOcxs2BweFg1dLEsaAkDTsHMtE+irlAGyjOEfqkZfNq1+Q8v81rmt/9j/AnvU/GeZ/h4HD0T2Ry
wluB57dH2vPqZqJcAr5oZjNZVhkovKLcxm2ViBA/cJ3hBF5zMxB4xpGXuFtSiCkoLhW25j5cKY3R
6BZeAWHZNxzWCdgcMzpEdtkj9kvgMoH29scNur9idPzgcx6cjlG40T7PkokpuQ+QTUw+c1CPXw6W
rHm4h83/LyDvn+h6z79qm+1cCG2GkcLLpQlV8vAF4CgnCssYyeD1zNMJsN161n5F0zM0tYpsplBO
4A9mgGfy0va4nUSP7O2CnHRIIq/ycrVrdNiSqM/+0O6tooEelRgMt2R9mcEKcnkChw5HJG2upb/Z
Qe4ktttOlLiiTFNsLZj2/8fita+sO/5csq+gB48woZZMHo4sxL7N1AYOfOxKzlJRSM98k2brJa33
BDQGnVZ7DfnLeufadHn+aaQqILeJasRhgtDj32pMdUOpmPaxX1TA5FIP27yW81KrT1K+IxQg/eTZ
7JqMoAr6qkeO4uhr+KF0GP1HD6bMyirzflQpa9HyO8sDzjLek6DogpsS4UD+WsqMFV0kozfAnqv5
Ra7ozxh4ZYeExjh5A3G7T2Um/+PCKExS3jFlkSV0k540jF2i9R0jXFOJZoyS6laicrKDlwXE7KKT
zWEYdzRt3k7UJ5u4h2skYlzBUjarNze0BDAfhrr1P1HPUkwTIHegeN4dFEmCaKaiyh2qlTWXB3CY
RA/XvcfeNPq9lMXyemPM6A1X0tReBb+NUPORCNcpAuHAhrCCqVJfWgb7m0bH7k4e/2j0MluIAo2N
DqPamGVkwP4ho2ERFw+YhNN4AkxLw97FirgVZJfMIfMauQXqtZjmd0zGI0njRyiBLjkKoCxFvV1S
mpWgFdor36bnCTZ/H/xaBPpmdY66OuinbPsUOD4rJ3fOLMpfypuYaHq4r55CcSPhpZ7OpO0XmIyx
KqDBBXWwp7HLtfWI5UiHJFW+cnCH0XbZrtNKOUP7IClFV1BXbCmKFJ8/B6Um3EYlLNNosGLxoDge
fUZNz2qkqR32jI1kmQ2A/PgXsFdlf38FZZzBKHt0ByNyOI2CkXaODBU2pYWw4AFDrrttPTxzT/Ok
bn70SfPVMAcMfHiIAmnie9x8xtXuh0qM6H8uGkaCWrMNpl6xXEfMlE1zni5qIhaaoEpljbSR6avs
ksJyG6uNQYfgU1FQJBZzRX+sxiXbz5mX9Yss8ia44KOKMqrm/2gi3lTEHaWEtTJVVD6toAGLU++o
L0Y/wDWuuSYZag1cFRpkh/vHihOxt7zcPOnXZpjB0SegosyddbFm+pcHmpCZr3uER84fre1N8h2W
d0gUjjJJlXt0Bp10JSFHsfm9duql3XsBvM/QalIEL2QIxfNGN8mbvuSlnNYSR7QNhJu72vjU1GPZ
A11tvAJtNaW9y8T4kN4hnBxGQfvaI2YVTitIlsmEiFEbbtUodpc/SvUur3A+p+yGKfyIA9JZPKVV
WpvxjDYCmhwmw0Nbz4dVp2FrjHogR/mHeDgJmBLGyIt5SeMNIHu7ky5KEIY872+/EIkbhgHw0dpD
xNdr7vHzmvJRL0Y1xHVyX/ZnW5IMFMCAlosXgtLOPfDyVz1VifCYLGz1IywG6f60zmm7MkswS3wW
7888q5ODyrvGUhNN1ySk5iDPGcXyS//BeKTZFZEUStoURQ9wt6VXaLr/QxolP7F7AGE0UZMXxt5I
LFqfuZphDiNe7iXBHUq8sBynx7DWTW2WxBq2WZV+q/lBmtl+BhtrjIVwtl78jnAfcz2LxR4tOcfy
ly8vBobAWMAGYhMQ2TfH5m1OIDHsD069PHWmbNCoMBR+lBU5kSvneOYO6w7hj81Legj2rEPJ/Ok7
4P7RpkDVW4BuKZBqfJX0g4hW3F5KE3lys3NhuDJFRD0tM0YEIcyNVmCE0rSYgjsy35fUp1yK3gbz
Dw7zUOUwuIoawOtgqEyrn1uFdiuc6+pDN2UTrspiCiUZxootWJmZUBQ4564qSB28DCaYVHzjym2M
2SGTqbfvYjVrFwaAfMQMXoJQh5J+OVJpxi9WWbbnp2m+SqH5qjHk/xqs2dbDLHBqeuXgkSC2ot7y
OjJsn3QAwGmJ9XKopA2DXHp1S+LEDUD/pz/eSKm0fRfsyDqebGt70OoZkVnyKmq5t+qZEduvildO
OhYupREQ1qzQ+uLTFPj+W6gIt4KmS9el/ZqcYjbKhM1lllYannivjMESboXS09anoG+M6wYMt3uk
1zzkFwKO1m3SMGZuOQD3bn6E9DlcxJ1Jn8XOdBFSL0JaUKR/MnoTXCwC23uUaW9qplzZhxLI4gST
MlLzRiZ/EvrLWskS+b+CrH/gs6TC0Y1Rp5VA0uaSsGBbLA0IPcYmS5xNWQ8pXyLYRWk2CbvEooyy
zsE6q24J+aF7NQxbNwlWJOV062YZt8Uy8CmgPSX1BOawbGv6EW3rbpPDT5dEZUeo+KZoADw8iaZx
/knF2EWD69UpcsW+dOdqZxlulI/hPH/Z/wm6703lXJNPNqazNe3h3YXLTBpsgCYbLFZqBPQegJId
Et/XikpTMnrLkQmnUdCYX4AQs8nS5ZBhZjOCN9QBhykkZpZs+l6tCEbsSgsWnsBZzze9A6Axo7jK
LI4i3M8yjDO9TcbStvh7hPgITOFZXZ2/VDy+yFg9G8hZY1jJsDmITBdr4aodn6/eNQ76IH3qroA1
UNtpiluenhRo39FYM5rPNW+GT3aZzxAkLK8ThjEo9v9E+H+/w6y2Vw5jRa2iBJYs1nFDqi4zRIdD
RuCWaL6li2ixQZ6XAgKJh46Zi95VoegVGfRDC4mJZRld2e3D7dVDHpyPGQ/c6OD19X3RQSm5Kx6F
wGJA+LEb/HHRvNu1zgqVmf+cRVJAuwZ7NSWmfk06A3kQqClUCgZ/TVr53sYByuq0/juUyhl1gwGr
dqbLa6n9DWNRlyR4wp0UOvO81PnMuBBsGBAXxEdcDaQTV5voDZsay/yFFxLrnSy8VO3h7MnCBY6R
cPlKGx/JXMYiTbna/D6dseFk0uJJuCIx3Vua2Gm8YNEXvbYsaXtR3nafuF+7dqrRzAkFt23qhgTB
C3+X+DuFmI5GgIvejdYNRHfixkqeGjQq7BldG5BxIRLc7JYem0x5DgZ3XqFoGvOteXCUMTm3gYIL
7NTxTsTos2sHx5J2h5lizcsKIUUaN17+FQjTNAEwUkF34vmXgyasiQRgYx7eQdyXrOPA905L1QSa
NlBP3AXztVUAP8X6ApXej/Sc34w9t5QEWUA7mEwlCSG4I5VueyFmL2Tu0+bwWS3FLMASUt5GdVms
40wPgIuZojptF8hncpnsN7J1NQlaO6pjNvsJLL8ZBax4PdPo2dRV/f1xazutll7zGooO7dRLAzs5
zMsK6LsaHzqKasTIXBLUtuXeLdjWCmW/5vmUpNhcWGB3kdTozcs1hlxADLmkXZ0feWcOjFf2MAY2
FkyOCZD63Xdlp2yBSYEefprl5Y/n5b866kkP3KOd68meIJXd9HcAkKgiC2qWhZs60HeqEkpP/g3p
cLMkcn0XvPPhj6WOFdjKmvCnmJCgsd+wtcuchPD8M3Z+smx0kMqsAEBfTrNayJ6lpXwI6DulgDXz
sI9gbTXuaiSSIF9mRruF/dhyt3sIJAxXPn9hRrH/NJbCashXOq6NzcYnaZdWHieRyS+E3ZKjjfTz
0j3NDN8IfPAgyVAAu0W1htAEnm+XtacPJl/ZiMFDmJDA0Fm/hnYlw+9qhjBEuSTn3M9JSR+0TPXj
QM7fyZpGniqNzxUo7s65/IyXS3pQhmDz48iXjHpoo1+RSId9THEE7BNvV2fmaiSeFyy231x+2VqI
Zi8Yhx4FEdmr1h8QWeMLZK7JIWmoQPr3fvoC+hEIlN4QTkIc0/LEqkZT4msCiXc1T5KHHJ6KkjWM
0ptbCnFTy3EigZpzdIG+dx6qmYTgwucMZgjw4VF5TPWRjHswlszfhsAa8JpioB4iPsTm3P/wVI2w
Hov45++ueyalnxE8dQytUnSXDcJI8UQAECOpiWQrm1l3mQtZ26RYCQ3bm2Ral5Tf/YXZfbZs0xU2
wZ2KWUZ9cUN/l+A8AGdZ6iy/dz5vumNs4czPVjbW7Dt3I1gZ2KeCqpV4/0EqBxzJ09/2bd3KEvtL
jRt2GRa5W/53NVFDxfsw2bTT5CKmU8imN+nA46iuCNZC2p50VdzKiwPsUcnbK5PjwjaXsGFsX2n2
Mtrtl5J+DhLUtDtqdzqZVtCler/zai9qStIX2pdEemirJg4J6T5BGqYRCDumSkcobbFkuGrSBomK
l6Pogu1fbruJoCaxMPxMXLtbHwYP9uXdHHKoXp0/7HPMmmcsy6xz3tw3BWXZEmoF44oNEuLRp8FR
3as8XO3iaDOgb3l06u+pr/1/9UbtXOzBtSoIeeYZ0xlKPqOzSID7yBVh46b7RrsBB5vv1Ft9QnxD
nE4X4+Ml7juU4xs/XamYoRz+MiZfWK4yVfQ1EQe54GdNR9q1Rid5z1zscri7liwkPnh8lMcs8OsT
EiVRLWnemi/xMti1lCE3yyqVCr2R9i8WCByJEghWY9Hlb6Zjd/dlk8Lv+a2VK+GmLxTtuKXsqgUG
8WQvwOPIkwykDo2MiI47H30iJTgwVFKLrOH4i+YYqBQ9xqZJgOC0d75FEFiT34PiLBz7nt/ix/T9
uR4gj7LBXOT1fOrYvVFJm3+7y5vaua8BtcdO/LQ6Irr52TaLlwKN30VhJg0vEPvh4I/h0TRA5Bvw
Zqdg2ZfeLRhQOq/JKhor2J7lXRmWN9LYIZ64ssMpr/z6ZKRw9IYx7ZlLC6DG6+aP8ah4HbvDw+dH
nBl6+0jpYraYsoKz7GEuiNHBp4swzuR/yUZxj1q3MIkkPsI6kIUQzjEckPs0Elp2/XEiSN5FZvTV
641lXqLJSH1IZ9hBbmUvRGoeOaBvq2+0p7TynW5SKEMDUlIxdsVBDQtWEOYqYmd+16p+pI9ZKFJF
VtgfN2wR4Qx/yXLBBsUsvAemE41fI86hBvT6b9O+aScqj8qP4SlmxMCdzeKwbqGsiR4EAy5bpxOJ
DlH9Z7nCiR+/FtaTkMl2FCR4tL9DxUwVzCNUgSJtmUMCoi47T1BrtQzE3nwoOHlna5zW+VDNu2r2
Y/ziDde7sOmd5yNw91hLSbHF4ymLGYQ1X041HkxlMzrgFsHvnS4TnCx7WFqP10fZm1yysmKbjcro
KWjgCeTinmq8h+efqfBVzJL7U4CZjlikCbDRcTCIZRHkYLheztenxjnVZqtmda6c+wyVNH8NKMHq
/YC1MBsEvxH6hXknY2vQOHKt8wQrOonwrBHRAHuDbNk9wT4xG39cVtwHisJEcvM3nG7jaSJ0USsy
Lv+FvJJYuqWE/E1K1D8kTiigxq3ovYJJWXiuaGO3wjgPW3x9EWoxhdMgRDv4FTDBiwwFZcZJFd9H
1/yCT/NY9lK6l1BympgbI2XgaU0/AvP1yRJhaSw+o2e3Vo+SE18i2TIQuiWMITJcP49LhyNyXxZN
z7Pp5vjH9hn+qx+ewnb+AEhIu4pH5h8qauxFF9b4naiQXU9lOv1Xa98UbOxtI+hgWNIdZnDVfV9Z
9J2eaNmTeFvpIsGwfo2IlL6RbE7tmrNuFC0rJDBwfKH8rhON3S7wfcJSp8SKs1JpW1oc4HinH9cT
zMTB+NnTupUuEaEfwWxSZaH/rjd9XlKWUWNuXcULLsvZ+mmw35ZmcLOdjgQKOJ76K9evBuxrGVfS
EbpDRE6O1BlwGC0rv+nCZfeiTYlqy+C3THxH4ZaKcz68eX8lHZ11K3IEVghZhIOdW6wSjYvX5KTo
VSvuX06rH5jUMAzLl8chvRBnNM0HlQQTkU0CRt7rn9Nn8N/bxjY5/ghq2jpLkFBlBJV5q2VZ8exR
4/ioFSSL27exgprDcIH+KJiS6EX/277RbvpnHOi+juvjyVnhPgt+LXV7DsGVcFW1GjqI+OmC6cZw
aza/XzS/n5X54LT68SxDoMZoEir0I1L4oB5Dcs4Cuhk90CL93j+L1UIl7Jf0CnIHbCFb4r/RarXQ
VJCycWKnV4+V+VpmXDuqEJgMktm2OAoJzEx5+nBLk7EizNb3eN2jxThQ0Q44G/ir+uWfZQ3Fom1x
UtLmkpLqi5Jz6aFdosV7PGtPgkQLdlBcC11neNpdlVoKdA4lmwyfeSbUU/N3Q9zjsfNaozh5S6ab
5dhCJCoxlE4F3zXooHmXkcwji4SPIjCKspiHxEyHr8pH+ZKYO5qQNGngcX5HfDzCNhb4QBgcuRE9
9S82qrlJHXfvuRhu8VvI1RVuMSeF8u0gVhN3AzrRj3K7sjcTcisWQhs+f3U9jxu/S5Cw0uL++r25
Of0AAjhX58H7LS/BreOmz5X1NpdDwVHbF5PwX5oNB6AVBYnaxVCx2sdb6H6dg3vik6yCWJJLmPVo
R6sD7kKQejMuTu2rWJL6mn1P1z6XahErAOsZWzG6KIIRi/YfYwictods+SUWrlYHicY0w2+aGXlg
7gLHC2YRi25lV9dI2WUJBpU/SnJ/JJHaewZpgfwNI5W2eYewt1tId1YLkUZ0B4eOT0ob2vuMg90Q
qTxzvmaHcZQ8ZO5ZiuIsmZWahJPwhBn+uSSzqGVeYrQ91RELdS0CyAhaaOtCjMH13qGe0AB/dNJl
diKbv2CLMbGjj3SsW2fbPlajmoDT9cgNv96dtsFaF2sqDtqKGKgCQ6HaQts7WmIa2FQ8JsmHFLGD
7fSF12Q8JnctKBojQw6baIKn83MGFSH4NMnzF+pC0Gzn0u7c0yyYu2ZiHKdG7S1FZcGr6HLi8/1Y
/vyKLH7rVkkneWUtVhzu2GkUDEt473WOXjEB8JZDvqIWLv8LlXx5MC68pgs5Q7/zx2lsgjd9IgeP
6v8MFSFLaev6Spb11yyRZULR6DZzVOvKVg+cSKxN4Qma5EWq5nUM3Fg97hAZLqchNk3UKu28KqUX
dp+g3jbGA6dSFVNNiawtBPd0jhEMavumDdj4cdNXwovzGlbE/aRuBW+3ehk1lV5ydxQaotrwcNNs
UKbktG8hd8pKwKzyBs3VyehHX9ShOxyN15xBzDJKhupQ3i6KIlhTQkUvXVhik7WqJopfvoLaIhH0
AQM2/1a3HvcnMH5io2uHchvCL2IwHshIe3j+r2SZVv9Vp0vcRMORRSvrt2nePKp8wJDJd2l4DnJd
J28u3jcmuEDkidccqrrLIgewsiE9e8+r+EdjgLuGv5V4x09KWNb0jXJiaZymGKXCQPYiWj73KhH8
SnATo7Q6kr/i6CW1UU4WJZQhielYJI1wRVmUaTUqQSFqlr8FnJxmof81nkzcgQCptjIMz9AyLy/j
WUIr/Lea1FlhjTHFc8+XMVwtozR2KS5wevglOi+Vjq8mP3Kqu08FyBWBR2HhdVUAW54EB8MO6+x/
4svz+qcuIaf8XXvR/IjYKQ0ndRZx2yn75A/HL03RCP8s3bL46D70KIImFTSZuBMKoxd3FGRgMeM6
ci+XPGmtBAvMFGbs4SSaktaBYWtPTuJ0InLG2odMm6qcTjr3YanSCZlARUTlaFD/wS42b2gkP2xx
aFoBx36N6D4KiUzhggNDrkDTlPZqZqMoBa7MraQzhfbLpxiv6wbD/lwg1bb2X/ChW2kqLXOV4fnQ
O2xfXJobsbzX/dc1aeLAgdQF+d5jYAOsrkGAkw6X3LG6YfZ+quT6wVVO4oHFBbga9t3YgeYxEg+y
jxuK2Onf1DaKZIM8sCgqO+v2cHvya2lU8JoaRVm/fLidSlmGyqb3+bBb3776F7AdsP5oA1FOAoaD
ZAf5PwQ0D2Gv9Cs7Os7WFLr0+3MwUbo0oPVj1qwpwjfWmyE0Ob7WuzBwWgcuhe5R6zQOnd+BzvTr
5nRQbe+Ugpll3w8NbqFQPeM31D+ekF53py2tDpIfxDqy3QNkVJjsnIOFYxGyAKvadU7GVI0J5jjf
z12L9zWYvvIQ1H10Ig6jCWazGxnZq1pPBTb1YxG3pknEWO7YcyxHCYxu2jwAmOlcn7Srq3y9Epf8
kG2JDd096tr62zwrKd1zGc080kzQ3hT95Z4BWawKOh3JOVmToT/qNUMV1/RNvkdb2/vUkLIPq/Gm
XLxOENySUhmBtm6wJp5WkXr3VOwV7cWG5JLTo4NmrlgidklqxY4P+rxGiDsY6my4+GZDTEQBot1E
8ngQMEtqdQAWRhRtELvBILQRED1GzxyGoDrVzWggrfdpYyI2PQ9wZeiZwQl6eZxp10RSi4TzD7cN
Xbxs9fgnSbFNNod49HXkJtmsnQw+1CQof31sU2Zq8Y51nrEIIv1E2IRoph/0gPiqBDvHQTaoUTWS
DvL4tLoj9IpFUC0+TSZNP2uGtMSTP4F/s5r0ysV+4Lb0k1EsBsQvZTQsbTFOs1qOtKi8I+tCkCHz
Tw3bhMAdEj0YBUd2jMSSm9SZHcyKGwU7m/ffWp5lRM54CeC2+nA/30H3/uRMA+TJqQw+jQsUsTId
QhjgHIR/5ogWYn70QlubhmfrYLdp9RpkK7fcB4P+YGf9inBsXDU2pg2zbMhA42mnejOCq9ccTeAL
u/WfEzQmy7EO97jpSXS8w7ZCBrwDe9JF+djJXOuHYsNn/zBuPRCj9Vv5t3w+QUrWmlh7jaYxVxw5
JVbEWxrFN+zdHrKU3siEPZGu6JFHmQmb7h9s00d6grBLzYCWLZu/RneY3adHCTA+dxF8n1oGCf4J
+ZY08QfM7ulvDiY19kwFOksy3tfyGbI0Fx6DyJG1V4kN77eRrSmJWS16nAWU0/MkqKuKn0iWYudd
yPmZpwEkXqR4sPBQ/MVqUlJctOM9nWoUL576orfLxl+gq2x9eLUlI8xWZCYhGjlGkF8Eb2aRqYHB
lfm3CJerhz8wZs3TqMyMzGhaGyfSSer7uLIrBpb4M2wIBAkSd4stF9XuKIuKfBdjT63dFx9FguLE
iAZeBsrXvIfmghYc9DBHIogsCjGQFIVlG+wxY+OJlMC87ye4WvF5JZyFgA8klSub2ig9bF2ECGqJ
8gmdDRV+tNB1wr0XzvnE2SIPQvRXK8nkgMB4MqJZYmFy2asmV2W4BszMKXOM+fI0MwPIpEFvGOnj
z4aMIrm0br8kIZCudT8jSWiH189WBBMi+Ad2XVgQ+14+3ml+iEoWSuZvI9hjhjCQKLtm43YCdhLz
MTEvDfBXKjwUeZ4dwKXYSOUDTZ+bG7IGAr0re8aXbl2IcxnZD7H3h6FzxBTsrMyhW4LfJQTyvmfZ
8D354Siy4l3SEivWnt2TWsHRNXwqMTVmc0C+7Y9/U9owsrOv1pu/7coMbhIyWvra9Iilxhc4Uvzg
hXGzbA5mnR8kMEd/1Aed4TzbXNenDaC83HOMUUAhBwh+XRltuQYvJXIHJYsDJq+UP5o3tM1o0gEs
9c+Y+mmAJ4d1duuHhbaCe8WNbVneHWrNvpblh31iP7Cy2vwmy+sMz2A5AiegPjN4GqpuT+ZGELTf
4ThxloSnUlpR22k9uf0TM7Jj6k2qJ/VzEqWlB7JK8AqokXI3JwbrTJddGzFb70530IBpKMWBpZon
0aLyJjH55IqjEEUN2+Bse56rOIasUyAO0vld9RWSVIdAGa4DhH+6K/2dKMm8Bt7Qwlde0TntFn6B
sl57nYDaolNq6s1szao/Xjy60q7Wgl5ZiOCZpBAqEDVspKCeEsFRNmpE6ScxV9q2mbqhroP+ytH2
BDW5rj3inHc/Co/Z24OKUaUtvPnLbS8KPFegojf+lq7Qga30iyWsihJ7U7ZZjxL5v6uP3XzdiX2f
t2kF0a9AapLZRn61JcL7RLbe/LY7L3vd6oXTwvFenXnqCo6euCQwykvDuMJDE/37d00yHnHUJ6DV
4Iij8nZX+nnXeTImkmWMzJT40qiVsHncdL8DMytAxd+HZZlee5viVvjCAJ5KOWl+W/iBtlP6iAHu
agl65gmHrsHa9v92mxGj3V63VcF9UI/efMwyRsa5+L2z4Pdq6wC8+Mitw4k3NCIfAlzcQn3oP4XI
07mf9Y/tTOrlTekQsptIshJbyNA5s/jqofpPdQPqJ1MNdY3RAyqzWOVa1YLTozX52vhhnziaDN8w
O+nIk3vgjy3aLBXj6P62zH+ONy6y6swV+0DfnqvmkF/+yFN6iH0M7J/4jMz3bftcmXMjdSvYhwHk
8Sqm2sy17ISHSdoQhfUHNM+fSvgRrKiYL7DNkGF9SG5kmmHwj4C6SJ9s3tIwiEBcLAkgoULXM4kA
vd4tI76trmTi5A4VuNdHd+gU0dsOfR0mwuSo2rp3g+1HSOZ2xH7cOU3fsSuApnR3bEwtBm133aVi
NSOcl4lGqecKzo9C4KI1CCrpEvijJot5Am3GUKqSxfddtSTlv07Rh6FM4bJ0KtU4Df/tLrc+fPiW
VXS1LrNSJ8sSbWJzuI3NEJpGj2AlfjHCVoeb9H7GdrXH1KxwWki2o3qxGNrfmPFHqTp//++fhg93
CHgPZYc/gmi6ZEQPxoqfx1Kskp5Rlz921L0kaf046rkgiux0VMj8Pv/X/aW9+QQksphxB7oZvWMe
5vH3SZx9KXuGLsPAGN5zSlTcIT4cRGhoueW5UB1xWuo/Rf+gs/WCfzcHyc89iwzfC9gMCt46TFh4
qi87Cn6jvFk/snd4qWxFv1E3gn3OCt4uUAmn7Sc0+FgMuFXQPqgZqKD9R3jNlqQjFhF4EBGn43OT
Y96HH8cjk2e4EJmskQFDa+mzxgwKdJYXG5qSdQHxhPIwc7yHaz6dact4OCv2t1Oyg0ke5xB+8kXa
FRjuDpjoDNysqlw4eLf3ovRyfnrWOSQS2wtcxdojS/oxtp8N2yitfFVDlPjoXIsBOa924nO6Tv/Z
t0wuRyQE09X8jjO3Ubr4EnTO+OctJIoeUgg5A/mbUjEZXeCTXWJ+f2ohYd/9bDGpJtLA/kt61JqY
vjOQbtCm/wrekLWYxHxb14MmOLz/vBMAkTqUmqmASF/IB6hHfs7DSjA6l054WA123vGii19O5x6I
96CK4paDJoyAHEZmYHw3eHTq8EipECAV2GeoQWJQSlvKQQNKeExaHMPIgWGOh83BiPn77Uk5Y3QC
tJpJjnRbuC8xg9oXEhHvrQUxKAyMwQqG1HPm5c1ted85ZmA+DMb73tcOBXo8EFF9gpOnfQupazjM
puxBMZIKHRHK925kvYBOFez8HQd6zmybgENSJmRNhQINokHeYW9zjMJvlR3afbLVqHzlroDi3GNf
HOJ6FANhwjrqEjFurk1YtSMfXScn/PlML5AwYigJ9iwVA69iAgkH0mk5HoICQrstVg+1VrsSYRjL
1WaO1b88dZtDp+baKit2Y5VVSFWcLQ1DNsyHO3AlSbqsOYQk1IXM/WOnNQu2dv9mkLIr4bW5PgJY
O5TIeQI8l1JQnoG+/4ikwrUTMu0Q0fxpEdResD42yJ9XIjqWHZYoSEVUfxJ67Cz7+7Pck1i8jGp6
jEKJMEPabXT8uOGWAiauQnO/k1Lr5tQvLcHq7e1Jbkqlp922PQPlXwI7YdVeVVCErOcbVFiIwUW0
HPmGUl4+WJAD15twB429CUiw6NgTTS0pi9ovLqOwSWl0YwfM1dpuQNR7RO2t9/VNmfSd1atTr/qt
MWsfAGVAslkgvWPiDCBQ1EnGOKlnSIcZXJtftABDjsrXQGeYCz0aqu1pyk2+8xi7YuidbDWxw0Nn
wP+pqZlh9J1AWi4BIMuenVYIpLnkS8F2/pS/O2puFBT7jnphW7g6e20zu2w/8HRjjUyuPJvx+eW/
yPtmKSYrY4stbifnShhO398OBzBeELWWrCrT8wEYtSYuzF+pQvQCHr8bGni8a/xtUsdyVnkhYUX3
jFy4VsEWK3mITqmmHlXys5BELzqMqHx491xnWvOMFvlSDBuJG/0y+HnsGx6gNga4nZxd7MJimr9f
mrRVIeCgZ5G0gNGuCkwNvMbLENOVYuGkDHW+07V9CfA/zhe1jegwellyfIQgdXe5zvKyUPygvBEN
p0sIBZdGxFCreZP04hTYdxokWZ26RNSnnP7tAJE+hV4kAHxlZXwg70ZnQvoudKEwjo+NPXKAquqv
JNQ7yNPiaPdexMOiIbylIUWyYojRNKze0sc4e07RAmuVgfmuyHhP4+tLB7j35LaLHXjJGjCVgDv1
UX1rYwRdaYYxIKUrBmmQRX8KXxnrhIReL2K3bSr0Lc9nhatFYSwK0KtFdhM9BzaT9s0xmKs0aYmi
WekzTwjoFdjXrVWCmc20ENT9HcROvhoHxXMnkSRfEuwCUKWoYX0B1vPW07Jd/KBumG608pY7pbus
O7ql8eC33N+0ItEXV8I8OiSaTaKA/50tZGqMSrckgYAxBpc91cfk2lmtXD/7ziqPk1sLhuZe0W9Y
HLg/0DWn4rA7ts5B242onJLN2xl18+2kyjTbaFIZA/SiHgvrWPRDXoE54Gs0sKD3X3v/l0Wrxwds
3U2+H2fLFcHFwivU1ww1tdFucEMVe4IvmjmnPsY+3XKMRaA0Ox5ZPD3y8lMcrZ4KfQmmczxz+4D7
ANFW3j5ubanBGpRrA3Cdnvl7MmjBGdl8iOMOyW9+5E4IOcO+GraqJUvEvfEzpXVXI2rIw2YOEj99
DfEthvmHxqh+cB8R+bxnbFH6jDOmcdRoCSZcwfii7sbGDkLByL4ZHHj2UGKN0oYxsnm84Yq7xxvT
w8XDigXznQC7SOC50EU5t1vc4U3Cd/aAE6KwSCLQv9isIfT27jJsdk+yuAvWQBXbsVEIdtgnzRgB
A1HVurP2h8jvU2Zj9yEY1kH2mqdhqKWlcfAAjgoR7fz4aoUZQdAqVLvARbzTfaoBWw1P+XpU5Usg
OOGy1lJfuhgM3neUqc+txFatezLbqLb6bzptkDZCOsrqcUa9hkLHuiP/ZZRXbvMYwEIWCdhwqrch
rmZEjMfvvuLo6DXDCXix7G7aVtFyCVUUkXmO+cIq0nz6nkLIKWY1WozOBXl0lEQBJ0MZIi5OGLgh
YO9MafVacXKdZ3njyC3sXVPYgBFvxQuMPx6WTQQpy1yHL6M4WYc5HPCj6zcqb/AHnvxKPNf6PSwa
ldxH1QI01glUzMf7H1HURs37w/+l57aPfJynoozvPB6SFKUrvHDXHzMO9N3CDab4xdBKEJwNTaok
ycy89QAdDM1kvviQK69ZUnUPZRNO/vh+IEnNH66rL0QRi+jgEJ5LHD/YiE+7pmcWCus2aKhXZeJ6
JmEIViHqAJCsOGYCiJKLMTfUWXaUwXrQQrYhBMQcEEwYAlTAF1d4IJ48CEKGRsgt6ZFzNAPPJg+J
sAt5HfcjvtckQlRTO0Inux1FNfLZlWq27OasmAwZp6GWreo+FnOKdhcB6N44bYS9WUz2OybBh9yd
VfNT0EfCPJVSWeEw9UHhMuMMKnX3wJmwiKTsvmSMIwCbCUxUmkL2IL+1o/WUaKVnW+/N2EEvewQU
RBG81TjmM4bUvltVuq2OlhOZhOPZycxAFLDbY5Cp7nqDAIdRLbUQAOTvkG3dMD+fTA7Tr/Kok4/V
Pb1d4UGvsjvuRmIrEUW7Y3wiB2k/wcgiBmlF6UA64B/DDKtBJzw52xZf0dglg1iFI3z0QJoKt9Yf
b+EfTzzDt/LZt9XKTtd4NhICtLCrYklinxicQsxY9Cc+NjZHmbnJXAx1mKl0tbmJEBZB3gfEBrwl
/UmtibxTGji7cZlL8k4RLJEezr+787p+couVlBms7xNjmypCFDKT5ocxOjqJsQ9VX2cfOs9U6+Gq
fHMTbmHuf2o90SBbSeHYzcKaTv4nYQLlDdU6Rh7lInFsgA3bXJZooJRzhpktkoA7nckBKtpmh2QK
2rAyTNWbNU5LHWquRku6+lDnlgb/TtN4HrrPZ+j/wR/8NgXaCIb8TNzI+bVVnFEFnoEi88Q4xKcD
mYS8bW9aUC/svqAbE4H6O+RnRwt836o+KfZcwTy+aDTyECyc3m0WD4ApC1EIh6XIh8Ymb78wo71g
2mpkof4spdEttcHM5bOepPMCjUtuxlxYbUEnGWKfTDCz+LZJkG+mwInvKfr7Wm4MGc9O7KgcyrBV
ApCORrNmSQ/WAOoljVOndVcS6d0Mj0LMiPxxNpzinVhgXVj28UzXIn6rwpNYtl5jmoYo1VaB0bat
YFKdxmI3zHyX/P1oGT1fHGNSj9W+Q+9xnuvULxO+rGbK4GUdL+IdCPamjwgwl6tJ7fEmjQ58pVuY
/d0rsl4szMAzLh00zPKluNICKjPLbkaoDh7vIZSogg8wFQuHR5xXEHP6Lrsykl+rNGSz/I4eQ7HN
61RoirJuCUOEK7sRfNfmtc73U2GV5D1Gg7m0nqKnUvS4+rQ6E9ULUPvAAvs1kipoAGp+nStENFRI
x3db3/9vl/iU6u6o2B/DtzXm9E0Xayy/XUC6+qNnZTy9g396GBGk2mTt8G0oJ/6eaZ0CRg8fZ30g
iwN1rjPMcqc/4rTuHECnQcGrdGtkDa+Ewks+e0uem4vcC4HfJVjUvkbVwG3L215TIzenwFZ6cqFy
2MtlPmv1c7Wh7c10yFDTWeU+4LoGnVYVVjwUpPaxGCIMk1SgBLblX0XnZOOBbGWmwhO0sM2WpCu+
Zf55QyJKkEgmAjHGklghZ5V5ZaKQpw4f0ki/9Ue+LxlB3ed2vfKrYb5bLJgnxdnKL1vXbYsztHj2
5gw5iFgRHJdfG0kW3Nf6uwdzDyXgKJQkyzPUeJ9xBwhJqzFcrUfaZJSCKCTBDUeklUxGRpA/8EIt
CP/yj7X9re7XNTjA2V7alAQK+QZEPjAtTB10qOWywGIM1P69xZgsr6MzSs/bMaKwW+aAXpGF5/S5
Cw9IhGjZW0wPoM1rkiMpL2Bu5Pxmo7CU6Pl6CKSgbBqgCbB5XG5Q/iQz5co/4p6LGjp37cSVP4ui
7MGS31QBEr7c5fEUx0rSgMfzMrR7x5ZCM0Yr7fL1Yg+dLFs3ovhM62lqVgrDhUsbLkAK61df3qKC
ITnEvEX/3hOskJRhLL86CZK7f1wddVoaiOMBxIzDQiq6/OZEYaIf/YF1QCn1A4oE1yRWv1ML4/1i
6hNMd1IzZc/LhVJcuGCir3R6DKtosr4g1YtgtY+QD2aMcRzzrTcWz4xpNkCEHEBSzO82ul0ILUTi
DzYT3y4sneHij0clD+sVKuNjgnuiqpTq8SGjbI3GkeYNmCrz0D5f+58M3qjAFEfhP8Ymgg6Sm6k+
rr+I/56NsPGsS1X+jg4QrEiPQ838rzZdRXexP8U5heTf9NVrX3bYMyDghEk/vnUrAflbHTSG5mf+
hkOBKxex87sebDQEMgwJ7FoRMitmJo6X8/uhimZWFQPPxw9+P+oyDKgmD4UIUM3H+3mmdoef/ksT
x9Q//dbuObxxzl5jbrWNMlT26IY/pwpriu/r75S0Cagd91CEcsDUGMnyH61ofsyRP6PHy7gBSH51
HDxjN1Req/xDmngka+jXfwgkr94fX/yZ7Qhap6W3BwK7zJN5dGoAj0cUknj4MIYoMj9XzG/FEqoT
dAwzaN9QoTJJzpzQZwF2jIB6iP+uC+Iux2+C/Q6Ys/sEBDHnhFVO7m775WRHIv4I7RmIy3dJWYV0
KKFmFPJO0VSxBiSVFDmgXeyxcghIDx2fm/4GnqcGS1Bk3bQzBPQQT8uSt9mq/yzaAL5NU2QdYAam
k/XIJHwbT9/aqmK7YUvW4c4g3XAwt3WJPppRIEJ6yW7u6iuOxzdfoVeQ/UYc/fqavRCWyyuNDLjM
7+gSl1LS7wBdGYMagF0So6Lkup1mYd20imjDvyMV7GvZHrtOx65+4TJ3BXTJQdiQzD8BomDnb2ka
dzUlSgPWzSJ79dMWySmBw6iRvsZvZkt416DiQIeglMzA860c7hZZRftjtglF1v72ouH7aIT16//O
nU7kcVNSSrlsJ+fS7JRW7UZ3zSYuEq3wf4D/tjg6vGfaV6KV6Se+6hNdAU44ijNotpBDTBTVY1by
UTAOxM4reeFknmpS2bvamPF7pN6bTWeGz7HsCdD1mkCMvq4Nl39775YxS6JzDxlsDeSB7RUcNo6t
TyWmAY/THWq5zDT9N0288U3CM8kSkEWdhl+JQ7eiSfGeLeOTVncrqGNr7E7XxcN/r6qbJ0o1GKFx
iX0yAyvj1k7JYkvD+wRljGuGE9Vyy6f8+3e9DZp9KLs8FsUOkNgQugB2sq90fzRfTWEtNGlTFRd6
yi2O2wrAYLjo5QYq9LeKiP3Zg+833oS3Hjwewrsm/GxVO+0pU7QJCj9zmKiVWtq05Ub9/5MEaoqo
JJeAcS2WnM2n8fdbLbJeH3vMkvZ6XC2I9iVyqzH9SfB4VLg5ys50H+88OqE0zSKBpN0qil8XMRv1
kTEbjXUj6QDebV1wLax7Mxxi4/FcR3vojBCRquahZsE+RYNQVgyOZ08iCsN43zaKyKQrVnvO89W3
Ye4LMQrWq5Dua7skwlX7l7XfXhpxRI6asW5iDiQqYcV9rucMCbMOmOpOltEErz+wnO01BgqvIK6q
W0iTel0V13QF8NSAgpBUehbWuQ0tc+3C/8N/rf1dcaZPx4peF/exxmqA/x+CWdjpZ7NNMX9ZrgEl
yBo37/46KwzAMX+X30YM1UpBBWhcEdRaTc5/t3F1jmR+62uOdr1gEbcIFa7968QS52T4Hi6E1wnX
aAztIeTVfRZlWGA2o9mdF6mwUjrdrIW5NzsYK3CDqPgYCfSLKVlk5r2KD1tq9bx2jRKIfgrXw3O+
XvgX1mkPBQ2TD392icZpt3CMp5vJg6l1dO3djbRtxL8jJDoKqRlokpsMHx6TS9rBRA4jCVyV2dsw
AGF3H111OOOe3Jp9nS3UFAzVxD4ymduN4hqh7mOfViiXA5GQ7AbIExrQnXUG/Hr6pSG1vx+L7r1O
neVt7slQ1IeHqAhEyo9lubMJqaFZ6CWtZFElux3DEmJD2UvMhIngz832uMgD7a13ChlRT3Tz+fs5
SxRqn/nNj+/tzAPv4glyqjDtY9aej3qTe9JyIHkdHtMZS93P0T4637Fez3mQD3d8tyEIODBVGh4m
75O4ycNjkwrlAiSA67hj9+ZNnHpxfEqlY57vGM2ZL4Hj5XamMIDRGlMeqRyBCfM+X1Yit1sYOfx7
zslu3IveGpDEPqpEDTbud8UbSYFgoD2xYHMbmxSsH9/jld+MhlKhWb+AgF0hXDln/EbfuKk78PcM
nd0g5HS6GhvskkR6E9HJUhCDHJBRiBrfrVqzPnkoib9V6eYZGrbrjVHoenqQpsjrX5rVyoDvPD7F
fL2Nr6qJfZSrdXKS6Okb3cCdozicRZwm/w4m+84j/9hHHxXW6OQNmPWU+OpDlCCQ8v1herw3ij3R
u7eUYvng3v/dUoFTgPktH7Q+0BNb2KhWsjwuZeUQ/mBN/8A0Q8er4pi8aEcy5FoEthouCNsC021d
2WAISHCt+0wPSRNnR6GzANIyWI83r1AsH9tfPWhcKBRUd6RXQuK23pxu7wOExw9l/ObRKGpkHoEQ
HD6zhXCbLUulcPYbVh3IA43i9hZQnK+B9avy3cAkRatX7iUkmnGq3qUxcpNo6ryG1+dK62Qrf4fQ
tNAob2EYAXHy5UVud/uzmOT/66NxzC4AwTP0/8IkAJEHWqb/1baWpjIRH9m6dgsmLFahPkBC87Qd
ha3vusMgdcQuSC02aEX1o8ueLb1c4SKkMk/HD3sp8sMavt4EorCaaLLTd3N52J5NUEWzDT368MVy
RZ5+ZJyQ/8dQySjVCU7hQ/wqxKD/GjuHcJM5hxvjtCkPWvF3P/mi3Bch8tgx/N6xUi50B5RBxAh9
SPUFbjQevJJfoGFSlBtRTEOYhWREXzMrlPI64U0gqmw6INg6z+mrJShXQ8TvJ0jL2hm7qP7qTfxS
ALLUL6NHwBBxrwYRAs64kzVJsRWANAKeaNRcYfmGQuX+Jyb6I3Exep6LZEeIeyYKF26XFJd3nkHn
/0mCkKcrTT6muMa5YTsU+a/lFDpsdVwaP6ThYSVjOhUNLrLqzTcEEKgkb8TC6U+FDFb6QAkoAbhS
xiWKif7Y/AQhacTA1OJ2y3b02yezwyXcBFT+aCR0ErFIh8ZAAt63jbxUTXpl/FbknjqmVH0tzA9U
52oen1Gn3plzbQJchKe/hKPbuEi2CfRTAprE6ZTaU1A/qSgf/f/DFdrG0RXPM4+Z3ulGMhdZuOdR
9/19LaTQrBp6b2Jebm5dseFUqpLVCENgF1/t/Ke8N6zzDGeEVDFyCqHz7LDp2Pyofdozq3GKL4Ne
CLiKq3FawZ3Pl9l0gj1krd0BlhzUigUVk/17rxDlMitfWGCEa3jHWJsR62l+RxlLWrDbt3SBbvpm
uyr0B0tvOKuwLmxaH8mUb1+WOCAagfWlpmpTyjZRlUrJIb7XFiMfUdV8UszXRMATBme2kShI1oIp
Lc1aylSFdb+l4IqtVe6bCYa2SUc9tXAL/TxbFXUEL28Eb9uAhXM/lC4iWADGu5EnNU73fZinoJ2a
RjC8kVm06TXf8BH3d64oyAwGmT3Sc6X7O8YCugVMi0ntgj7D+tUuH5SC4NvEMtgmKtmvGU+9ia9e
FiAUhoI0cx0hSxS/yUNNEHL5rdaqCN51KIhi7XMiHRutBSnTO+sTFV/lBhTcm/uIjohsDduR+teM
YeKBkjmHKYyXZbuflyDp0875UtXjonwF55walCeA3K71YI++mRvAcOhe8LBkOgM3ZpFa++31TiVt
1QiGx9elq8a7pOZZz07uDKLgDwfT/4Ugta2fOnXtA9h3bQEsAPuzPa2XOsUju6cWekGT9Gdcu1dR
6HQZD+r2IiUVDMzLuSlC624gBR2P5Lr/We7VIud4HPZJH9rQF5URANSIKhk8GF+oj5rYtQkUckBz
6JcQd+fPDUfOALqJV7PLSt77PfX0M5O6DTnDwZ91RO/UGh632wJvoCk0QLJsY0IctNVeAM/H/X5n
WvFY7wPLZbhq0hS4WL66qS3+/BBvDnHmsG+gs3mcLhLknoP+v6v3Rp3ErQ/B0yXx1FaEedUvq1u9
LmEEKFl1UqRhtJZpRzgPXUMe03RzeHEllk3B2wKqXys0XjW+ziW271+iB8B+4uC/ER9XVMjYIgiQ
VOuxRP0shYrGwLnDAYHp+fEdM0wKDbr3Nnlqwt65YijxuYkgCClKOe0gPyW2S+xVzgDQcpC/bvRG
RYA4OKMD4DjTxQwAB+whx1QpBrMswZaaXVpa9uOVTd4GxrDJwtEk5FtH2cQAQ+F8Yv6IIBpgmdUT
OTZOozqMyLz7DLNsIshxPu61WW7+rRsK+BXjJEq6x5stT5DHq/6zc7uFDgZd/fBmERXUM8dG7fJE
FPX9K8ugqSt19YFRFPKgBrjEXlZeeMgcQ0aCa+D/dpUuE3WCcF8vN60Ii4DOSlJUyh6NwO40dhEA
8kiaT7wy++q78K6lPpt4HrezYo13Y2GQNsUDtWNJmLtDVAW833OQKeXcQDaNfCkDCKW7TMZUlrGx
JB76v8ZlZcHzSdWW3H9hb6tsnzljKr8XB2MSknY0eqGNi+geNJJbUDLeIHZNv4YFrWcMZgC5CRLZ
3giGDS6lsb8dVb6bJ7UOfh+wt9cPwsGjpW3yV+XYiXVtDvEh3bWOKQeTnSJKU8Cl7SPTfvyTj1sN
DCTRzYFSUHjzDWOpKqG0HnZ1BXm2ymRhfe7CiZzxu58WGKSbP0HWQJm1NcqV21G/eo8UE/GXRfwu
t/V+UN2pHIab0oG5qv56Z+S2JkxbkpebM/Q5J99VFAGokct67pOj0RmK3l4ZS+94l+VlNYTvzt/r
975T9KrE6Buqv9cEjlyQNRb5vRsPWZx72wRwJyaq+A5cEDIl8bKccpZvQNjTX6SLopylw1IuQDCb
Wug3LzQGVOhFLttoYkO0nhj7o+rpk4SoTFT5k7US9zz1cX0ps2DYDMVs3U0+aXgxSo+inaOly/Oj
s8sI8IWAczS7X9Nbn4AaClu0vBRIvKpNTXXM2UF9WVBP5hNVYfMVJUH0aADcLaz0H/eCyOaDiwRX
AtWIl0kE5aWaMVJIAD92sXUrSvdmJ9HlupHtWjPj4Ej1XjxrC1P4McDR5s1IY/92O23kpz0MfkXQ
TrVJwWfdNCDvKNQMXjfiXhpzmWIkZ+w459JFVbBHgqeD/3lu5WwkKdyXDluNosTSsGODt3BFrwkc
E/rAYgwwd77tNiovoz8SX+Q3nJXcGywostqINGUo3wQJSBSh+A+achBKRcPU8EHMgeqQQtlQyKtk
FHT6xL5SwGSbmr6WEXDW0+NzXDe2n/P48LMb0ik2zSJp/EfN5jgkqBQaBm1PXxnD2E26XiHQZ9rE
JnObKmfaH/kkpgjtd+Cvj4XNM0C/uC+ofu3oWptbF8YPua4xmE/jQ6ucDqR76klIJH0XdeSgwLUa
JuefjtEKN+44j2bgmEMo1F1dNNC5c/QZhdKTwFd3c7zyD4qu3dRemzPuvCG7PxTC6dt0QdcHbZsX
4OcHoY8FribJLEHqcwljW4longx8cbBSmsdq4oaH8e2ZzRgcayvcftNjAPWEUtsy6o+nQFPQH89w
XU9Qlx/0PKgIICIBvmw3g4cu24NZv4ZRae/u206vb7L7QLoyuAnLXjInQI5CEIZpjO+JWiu0CfRr
+yMMfam4RfpbCl51DF6NCQCEpPXHgAhnYQz4lJ2VFZ3RrRFjNuin+gnKm3pxhYcBsG6gHmhjZq/J
siB0Ukd4f+ZPFpn6xBf3jx+c2GOVAhVPI29wGQ/3Vj7DCmo6c/Pv9PcVIO35njt6RK+hWU3stG5n
TXPvfeGyBcImCzkkMTwrzWQJFJoQqnpZc2t6PqmPRSLUMoQucq0hK+BlIUGGxmfRlPPtciKlB8jj
PQNAeMv1UtNfAMVqyWV/4P7pV3E6Fxw+dbBHEnhOsHIhSEOHnEoJ3j4Ajp90MaieOHr9VmJSBN2h
3svU/Oy2qptZ8/3pfInEGRrxEmzhLptrAExPZLniqQs+xkbjGNW3YRw8HgmnffUWHZWq43eox8zN
O++rS0tA9DVg36JHUhIQmBwVpotIkSXIQUoDGuR7Xrq35JVi/LYnbKpXRRNHgSJJh5t5CoZ9Cj8z
UMbSseFZl0GxRzlGc8PyoyEX3CwYmzskNfv+ymQ9RYeOD+v6/5f3t7hvxyMt76MyQjr61nc+YDVR
tBRUE3UTAmL3WX7fwWbhnFUGSatqsRVi6AQp4iKBWTcFmPCbCbFrXjGonUJfVod1a2N8CIVGohag
XatXPe6JgqZ/HM8sNH28rB/LaoQ0ftmufhmRYMmsQ25+zTD1z8Zn/qOaGysqSv+9Pi04yOz7pGiq
NFTFERyaIKVFZ3PxIv+zJpIkZHVPLeINSM0AIZUEhByvyQ9sMUqxjp+Trifz6Bq8J4mPQjX0edxQ
ONqQun6vsTDvypdnVDb05gWQE3P/WCv9Nx3JxeorN2gSJPPtsfSxripDmbUFkFYmcNLo2ATc8DxB
xMBte1zeBVwuzAmfaKnZbHCYgx7HLHaguVEBQzD/XXQCXnJQ7cFSEl3f/PAmcdVeti28E/6Bd7Rr
UkaC0CEB2PYLnzBYmlwBRxG2HgU/Q24I1Q8eBUHQdB8EcLl4XKjfGi00Rfy6rI9kn+OrRqklrAeC
uClPMLekznRrqMRAGeaeH5Jp7c2zCzSEHjojzLjb/FCZuIpgZvamn7hkM6rVUgVmrRfwsaXqWWv7
nF7bcZK+FWZOQ4dN1A3nqebzZyURLBzrADvt998xBTwSeXLJcSNG57MTwKDbc8GncJJ6S9lPhunP
/zUXqqart3wNZvcxcWXkzDPw6Ur/mwaZKG5dyRG2h8mad65A9msoyKozHDymurCNCgp2XKuqPfvd
eJ4XP4p8JZj9F4KNChjDA4UvVCKkXxdyh+41N4H4BemXkvh6Bf1rElFiy9OPrJbMlz1yAgOPZ2Mh
JEoDh7sbk/uQQCJPmUkpHXaPJFQohTvfjbeHj4SfPeaDNdt+P860O3N2hbiB57LTrt93r01R3KRV
44AZghQb5HfRlo6C5KuW044xzt0FlItaEG7a3CJUQI1MJE0qwTx9QzIed6SiI+AqkBwA8awb6a8A
e/RYfY8vIWqa+RwKNZuKQyOfh+A7C1oqcmnJjsGO+QnM2Dd5tUtR2H5qvetquS3gFnEW7/Tz/+m0
udWAz5siKyuoe9JZ3YJrQdWxgSok++YTREvsSXU71ioYNbTJThj0alu9IIbfXvbOwe/P2dBe50T4
H2Z7iVgnRqN2J0lyiJtVb2W3rwz2KYaP1b3qWWm2XOUVYt/u7hQSVuKPihZzUkKvEi5RMOZ/KhfL
Fyb8wwYvRdbuxY8jaRjEL3qKsnoIeDSB1P60gRjej9cM66t1iIGnMHzrIJjJoczhyojUSakFmzXG
JtRCwq/GU5MM/Zhs6DYvRie8xLP0+NB0NFUgfZrQzFnfk+lH3yCnDmwUoAl/YrJi/NudR5NACGrK
iR6S+6ab9J/YNE60/Fe2CkGsFOhQBUsiHW1q7zBOpGQNVnz/yr6mUPQA11Z89sZ6A2H7zuvy1nsE
vbzklQMKvMarBozFwsfq0ecL/TNQDv80HhSThGHgGjnFUIBNzIvrvE8Tp/uxDobnOf0AsIusjz29
N1PTQfs5WdheQQyn7QNvMVY9yP7A4sSb0l1wWodHn/hPcfxUzAwaT5MiwX41+KanNsNNE3wftlQf
ZPBjdvAe/YBt07UodpLfPM2cF5TvfnPTMOkXc4hKTKFcYkKk34AERA1SghlTpYNGob7gMSfFeb9U
WPFASa0c2QR0z5gRpPJc3JVkXPFy8j82DscwuebS8Rxf/tgjszutbo1F54H4eZcbzGos04evIW6b
qSTXsIKExAvBvd1XQelG29j5ioFmdsLilLKBVWGKRnfTg50ghGUWgJmsRJ5jpymHhjSlnlcsqRoN
s8ECH8JxKPVnSwMJZIIZrSTQYXb4RKCpquQpA/2dnkN1QqQi/7x9RWAGPVOfAnAmjYM057a6+Wni
oOluHTwkksWQMkqVhQ/sYKmu19uvVEQtUEbbsBN00B2ynKPOblB5w8jBVgZxb60E3Ag8XilnvOdf
iI6QuLTUpQxUOs3+zWRpPl00Sm2UEIx/XQuIjqOKc97JRx7NXaJOmRzdsqJhEt02P1JXxXoFIQzY
zwZexQRAxT6C2nPn1W2HdLdUF4Q1glXs/LUMuzbgF/RrU3MDmz7D7jG2zN5ujKdOJnvdu4z35ohl
ItGxGctRToQlVZojN54+AkCZpMs3dfe3/uCaviMpObILyU8CuQaNRmv8ZVRt3LhUDz6tXjAE5UVC
wDtvc9WzLeAmy3HCuwyiiAvY/wpQRWHjzZshC8uQSdco8okfYY3w2b9D6FUcuHASHC1/POrJjJJO
3SaXBE4a5BPw9uxXDZe6ODPUnvvq49PCKe1a3JIDvy29ZIdIcLmyJYsEqbTtKcrxLI/cB4HyLgyq
XxmdQjQldzfUcZJT8ddjm1GIBqR0XzL8Q55eH/0sordIx15jZbcFcP/KYBaH4e6COS4hfuGKe0Fv
4AWYJhNQtIfpUsmVas9jzWRLxu5aEFg9nUsiCJgydce/fn3m3nznM5eE9qP894jAqdnBgKteCMJT
A7WfxLGkfFJnX/AEByhCBZob5YXgYuZPw0McYAf3tIt/UaWiHnr4GwbfGQDFG8TkBDDYAi25EVlY
LVrwC/Bn9SsQdmL9wBGPJRR9ChKhBvJt270mkOWnS4a1QsmV/3UOKCjQH7IT2hX9AqbIUVdZ+n/D
We9bIdbmyg0WW+7mLxo4ofoI9D0ws9KtH/urnaYF2JGUOyLAllz3N8EuuuzKStAFENKjfG92fo+T
mulX+lrXCCEEY7spKTzRBDCXApEgYhFsSAbwjORE+FQQ+NNIbm/qHlyK76DYwzeTKVKMA20okeYR
F1O5B8GfBs2CctRaDxVDRaou+I2muWd2J2E9FHfmiOnR3Og2vyKDcJDkNb+qRwlKrGj12Ju3/jcu
VZrJveFK5LzpPrXvkIikzQ/wZk7Sun+Lus4D9i/7mF4IKSVmkmthGpkFVNzwtcJlsYoDppfDtQuc
isMjLdkBfI2hIbjlK5FWz/bXMNzXCQjCtAI/0XLA9yWp3wGhFkta1aKBXXGnaRcZmbkjUXlv0QO/
50ZpSzD8JdTGOrDOWDNeu7lyBRrU/UA/J0CsbAVvGeFfmNewJ7WVt/R/n01IIpIn3/cPBIJ9Sn6n
xWioIgsiYWQDhe+uluwClGlXm5vf9K/LC2lnm0WAArpOzMVZSyVeaB3EJIH6XoiyeoVOmr98beHg
iq5jHx87JCfXHqfGyRm1BQp8PJFQ/6Atqfpq4pHNOVQDMpSRSzJ7bUEgqCzitlrmO3TBvxvYN1e6
yFW/oj9hMRudzfsrfCLYMTYGpQxEVG1aM/Y9hofiJMHop3LjKKsr2kkwKiXRrwdjo7OvyAIh8Ks6
fwr9tSz9uBOQhrKE+JjDkP8NfE8PJY/EH3ja6py7ObddKwbbXQoEgiCwWpeKoFvSvDmLTC24XklS
2hNaSyS4/aatgdjPMPkuJKIeDfZhdwcF/isOPtQ+jdG3CMzOhLoSc51S7oAyjUbB4sFpclrG1hJB
/VsnsK58H3I3k/v7ysacmRd2lUwXaaVXZz/J2dZnk41lKfW/MlbJJUvRySryHKAJinL6D4AScbaI
lUker82IgvdcS63m7KuP6djsBDp729PmR243+gzSF+hDozi4ddGsqdN0g5uzCp1V+gerowW8T0lO
45tpAhyGcN0qfzQpUQnOPv29kNnDzA8lUVezlguOF+gv2E6y2yb0vSb7qQwl5R+4W557m3SAmzbQ
mzTmCPEsK1lkerXakMj1r95zAL8MQUGpZ8XpY9o+yylV6pm973xisttFixl1a5kapHArDi4qM7wD
Tp7lytKenIDCrrRrWXmz6fQUvbhsbh7L0udKC6aflC5v/+OWwcWGsqfailW2dUENXsTnPqdKSqnX
epGmaNobelOu0P8wn1HxqBoZPr+rU0gx7cdlGsHVBh63CcsP9pxcYBiJ+PbBT377G+KHJo9Yrlps
D4QMk/JAHm6kEwkNAd5wO3tCU12T9wN5xmR/5dg7SNGI327nm6nByT38R9F9zHJ4ViXZfCff3Ff9
bDkhzDUDBHeZ0PkNczBy08FQkur+MpEKRH6CKoKMTUKzggERN3RemZnNne6FREj7JRQn+cJuZLDa
KZ6VvTfMnFW6vwru03Foi+9YME/C5J7uTR0rjxQ/t7OXuBABOD/SpB53j+U/B5hC6XvN96/iH3o1
Ouc7PtxDOsaIU+4CO+xMQYC6Xz7StCFonMYeYfwMFUA5MAyHcg6bmbUKOfogD7s3UZquH/hRNs/N
PAGHyPcjDxhG1VAcx40TifvLtBe+yzUu8GhR2ATOSPgOvPkhOUXifI3XslTyYkl1oKwv6avH8eys
knbna++KBxV9hLF9h8TqnBupfyFSLtnJptBUNMNk40LbrKagIdGhQ/zdkBmuZSroIHHZnEXitYED
x7dHl5uCpKPmBclwb9jPCXbLhrvTIAbvrm+BxkF+KUvDoIFoi/e1QqbTkGW/78qRIpjk/sumDpPL
PMcLpsHto7zb4jXtc7YQhlMhC6Nc09ieoOFfkHvrVTB5VEsu6H5DxUneOLJq/zkut40OYAHwW1gX
YYdyAf9IykoOn83pdBmMfaN2kcnWbC9Zxp580RCv4FkewR+GDgGNpsYkXivPdTqS1RV+e3ncFWy4
iMe83END6TkrNPhkWeb6bXAAcFGvWTatkvQOh07na3eQZ3cPpgFDURRV8+AUIGayw6LccUrfv2Lx
mOEOmKsIPPF6x+wsx/P8W7C90kINg57+xIqPJ5qYyfyEwgiEerLS/S9yqEkxlwYcZFTSlRK13kck
fm2mMBdxhI90d686ebceKwpBOiZn/oyKsVtzAs7yL3wCEdcJQtFQARcl3d0ofFOKNCqx9jEYHmg9
fPRpLhz/XLZPNRrX/gzBbFkvxvVSbK57+DRPjEdFYDMW2Sf0NgjLr7wDRZt+PhRp181NtHn6aoTs
JrkHsZTTA4NpI9pkY+zw990MflJ7WuFttCidg14pll0l9tO/zhYKDtuFWT2xJnUO7Sp2jART3uqN
cA+k1kJBImKaIZxNxyj9N0v/kmi/Kt1FiLjOFMc6W2uz2+wMQRzytit5uMNG3QgG5YhaTz7KtxK+
cwSJi2QMWa3m/XMBvmCTam/BYSMyvPSF782OgpJwgWZFbvI4TT1pKOpz5Ws2u2FVwEOL54cU4Bvi
BpZFDqySROFYDpjR3hV7NdAMC6ZH25hR91IWYNzi8N9r1/33T7TCVtNe0usoI+2YqHQTEytKyx9q
9iALgx5dAmcux7stsHx+LwNUcobowFUAYKoqHt68NsTgTIPxX1aDmuTtpDxCI59f7ibpwzm8Vove
e0RHyIxc5PMH5OiqplxiMahs54NgtGBjLtQbkOCI+GuCbyXfMdOVcixxkaqNDG1JZ1ERU01RpVFs
Xy6wA8/YJ7BQG8x3YExRcY0kDGKmiOJftvrbzYUKHIYtuG8Zunzb9zN2oDK1p2v/c1O9bJRMspD6
qS8Gbi8Oc/47JiD2/q0/6d7Nadfeh9vTXN2U+Ffj9ZeYaMIutodZsIUHajXTKa+A9bfIa52wxdBk
+pzYTAdQUWH1P7Fww3l6/VMpTf2Z584CML8ioiutS1VpXHb11JC3Dy7rvHSGDpasDEMnkwhvdrgb
DaXSZC7Y5Tk/UBItF4Z0X2HjpFEWOGC1ic2XDjio8wf+7+1dRZsj0ME0ACalM4HlPV6VrPBasMaA
tq7aN5zaDqO7MYFTZnReIJO8qGQ/nmiZqwUFMd56nxakwnbsKUMyBengJjSQfgWMdmLI4Ln+Hmyc
xo1hyGvlFDlO6JJEMn70ep4gu7uk0g9UBPLsGaqm9GB1K9uHdmF0SgAN70KFbfYtvxXDmwU+lg4I
+baVawJuj4F/puDoSaWn3BJcy7mHQig0Ow25rKvsX4dKnokHPWVJTHXdxk6+5cEdVaca7cOwJUj2
LvbxwN8s3PG5XD+MfALZaIQlILpJxZlNARaAzRslzUy/5wwZOxP7Pq56YWuYNvo2H/bzUCPdxi63
hKa/VC8i6nM1w7gNeYd5IifaK9ghpdwVVROxfCFEMfXZzo8vQ4DVKFR6Wfvse/CxFomDAbrWU8Sm
nkq8WYFUQZl6zUxgj7Rb+h+cddinL8IL2rzFIsL6h9NA+dvN2EzZeI6IRo5PmCSYksIsbsrFmdu9
YZakDu3b/qPcSt2MUqcYDHgwfO+EIB/hikrNY4pG7vrI/7hP3eNbNgp1iofed761qu0kzMB7egnA
eRGE0nl9y0BS/E8M0ARNbvZIwBdnkYVm3hZHnekFJjP28q+tNaupx/HxXDFjiRVssgQy8cKQAlXl
W4eV7XO3oGDQpLdOGp7xnYEEGeGIN/wbH2oIoDmPXWM4iFqSOLDu7xQsHCG0tsqWcuBCNF6gA/5J
ghHSYFNeCFOL7qBOBRsSCBjATpLFJlTFKR6IIKiSEUJUMw98lwe6vlTxP3W6dDx+UQCBywWc1Py9
2EgxHC/Or1iORrzPMXKVpcehUOZBD2VDJAa2s/3lK2xRWpVfhRP5jsL9ocYD9eS6S1+oJgsPTYvn
kjAwSRYsbNARDDPZdAiGUrCQtOKk3RoH4exHJudQe3eT8kvMQ1TjOejqRee64n0kY/HLmhPKAG6t
422RwDZkLPjoIS46CD6BQQNuHLcZtV2TuH41H5AUodBVjQPSVUbwdjA2SEaaBqJ9ayLbejstzg0b
YDYsVlHb2DSYIe23tdxsDNPXAdHBzPylPZhSwKrK/tUILqHwqDs0MFaz2I8QXt0rdDn11c7CV3AI
q2FRVZPYymsJ0XwOO6Rp4g6MwTXXSDE7EG0HOpY9icG7cCYqTM5c2hNEvs6SuJAQRhFWcTx0cCmW
U6BvNlp7xVIKT8f6AIl9aCJO1GoUmaufZbo4z3DbSHGv8cj7uV6ryoBNYm3uBPkFa1xaE75gspIl
TmL4NiR2dMqxJ6aagtIt5x+XdBll5EwKXJD7O1+lsGTVn7JaLumo6n/TUrsTev33HtN1x9ZsEIdO
f+5obBVoPEOGkz2+RbNOdsZaVd9JzBTxesRyORk05dpdvxSkIcfxWQhj/GUFP2uR9uQh7jplFTui
kcUpRXuku6GoU1Q4kZ55cO8qe7trDeFXrYnSr47qJjVQ5qkBWJ34vFTGLsoGg7PlV9IEGERXjFxu
VsMSKmvwIJUi1CH8Ia0ClOFeoPPEEtXyenFY/0a1p1uMoaEg2t1ryCNQOe1jCxL4k9f5TZrkmfTh
pO7FyOwzv4vCqZp1dkor1/OxLCwurIYJX4cyuGtl7QXyMrBwCyO0gYGGGIBuIC68m31lZaYqKkTy
OJzplzIfGSsm/5p71CDPuUsS0XbaXBs5iJz3ZOACX44XHMRTTFPk0i3qNvYdHOCptL7JWTrF3Ppi
XedTsFbLYfg68Q6EE+m2JF1x+UlZ2w+set5qkpaouMWlxnfMypvXxF9WiKTOztl4QbXEJBxJcxD1
lJnNNdmaY6OMzvCE8KwuKwjihXWsDxvu2hbKFC4hmGqkg1aCzcD3rC6sbxRAxbE1eIq7THiJxbQM
lMhfyhvKC3sE4He1iwjEsXTJTyplVrUvVwZX+sZoD1KGOHFmt4131k+dlkMxOLoEhJAlFTZaf9QX
Q3BG65LFJZ7CT3+nt6CF/hWes76EYh5A3Fe7lzfBEAHM/lES+eqUxKBmc7UGlwZZBtlah6yPThIc
o2FH5yF0GXHZldhyVuLZqxWZbxBcOOqJN/V8/U3rScs59CvIsCRkpCBxkOHyqtaElYmv9vTd089y
yW36zmdE+01NVj/at6dHAHQRX39H6iwW11ULduS1MWvRFlBetSP57fdTpWu72Inz9fXjJxAJXDe1
2Tzr66C/FdYyxeVFBciq0HoT/RFu/KKY7MVWqDrdjUx7Xqm4EpzfWFM9Geh1Ejjr6p47mQhXiUn2
BUKcmY/mj2xxEeZQRp922sDdFWrsq+b4rAA9GCwA6pr3X4PHEpc7Mbp+nTpHKknddYPO/cFseFA1
IVYvgT9HhLffaC+NFXw2tkvxFW5k2QrKjym1+ui4YINjjRMjblxhf3VcfPjo+jtuB0gC6fTLrVcA
0MGM3zsjqG/p4iK+mLv7QA0MHZjRiEUr58Uv3pNkNNShKblH+nzvbf3eA7RyfFb9/pFrs/EQTcXP
qdbZVRAJ2JmHWUmUTEPpV2fXiZt0sYvUgL/4QRLoemvmZTImkceM8PQf4DExTTS+Na+QWITcsAUT
sAb1qSsdLt2rDlNrpzzf6zHZK219rLmhN1uBkIKR/ZX7FJ3poUXNairjJt3WhgsdKDvb6ZILfTUF
hrZS466f9icInrBwizRwoHOZ+HG54sOzpGoeEqk4QubzYiQ9bDTQ8XFA3dOspd13i48Q6Rju551a
6Ye+5F3dfcKkZl9OFQXSbtA4GY9LBD20VCvHec05DQgA/3jKliL3uqooLWjyVeZbUiDO11KLmehJ
MEAmzDsQdE//6gq+p+nYKiegfA/ZX/ArKH49Fo8IYd2/eIhJ7qXKZiyf+2GHomN+25m59eVi7Xnl
YTtg7yZiNg3+oGKUMSKFI4TaMxW67aEjgAVphzp3ZqS4611+JsFUXIxh03U20JISUbgyv7VOLhi6
AQjG4GOsHWv+5GVX7Mt5N/D61lOeNUoQpVoP7ypJx0gW+sNG9Y9R9dCtFbFtERU1Rh6UTE7+lhv7
N+mqzOtov6KjEc4zTOqH4vt7X0b5C0y9OvbQJ4vY418mC/O27qhKAICh9hLwLE3rV0n5JNFaOeCP
O8ZaVuLNrBUvQ+a515YMI7pIIiZwAWTfwdW/wfDmGIVR65rmyKidOnPF5Eg6VAguu0C2q1lsST/s
jUvR44RSer4hU4ycjc5L6ifv4H1YuERJ00hMKQdjRVri1W1ZxfLTtQpnR7eYwGlrT1oIfSfpIzIF
s64YhgcJlZQzxA3YiMJsT56byZqO9Fdk1QJZpnCEsDPi5CCJ+EcSzCR0sqPXdYQS1wqMt0HKfk8t
i/zZNOGJw7lhXw4a2vigP4ddg0H4KLuyE4BbtydLfimAvXgSuUZi8Un2bhhQU7xIZlu9esqVYEKc
eYqjZZPt8NTBqb2yeHBnJGJ/AjToEbKZNoHYBhte1gA3lZ4er0AnJuGtgiL1E/0H7BP1+SdIWNBH
C5oiBRIyhHnCScQbWGLyIUtiFm3IuDPeriFNC9olGXq0GMwMsjHFw8tSsbY28NgrqT0f20nm28WJ
ootZ+7aCKrW0+6nfFFhcrzuUECcEjfN7zRZkwd6OkI8GiKP46myrw97ai2s5qRl6uRS33GlI4olN
ie7RMwvdqsIjkOC4ootSGwJxevQnmlhu/7NG7ve6PBCDU/psW9oFIPBczFrcVgk0u4rNdiWy48T1
lQZZBXMW2ikVQejFZyqi+QoCGksfRDV9VarfpYVQbePf8lz/F+HJp5C7rV5O20tUvxn5iVU3wsL+
soURQ16MqYht9v+8xpmViMo0/ZC56e0DN7oHjG5O1rWXhk4rsO4ud/SKurSgAxF6cJuYeUn3SDKQ
J7ImuqVV8AyGxCTpnTB2I7cspaeAPdDEWP8GspxYXf70awdlgZtkyWh0knvbcDJObZ2wgvh0Usbj
Zhev0oYqf5TvT4uZwJmsWvVjidry40ZgH4XqeAUZjCWlRqAc0Kw7Yp567m+PQjbw5eWXphs9fmJC
6YMfCHFp+HVtgpKs9fIRsND16HrhCi6ihRgbm5k7FyHIucV4wTKZh+Y8Fzp7SPkUTxjVEc0/DVtg
H7KLpezFanpyZ/VZ1w7zO3+WnhMCJ0QfvUwvHpYxeX3RBda0EmWL/KKF+K+3ucDkH7obyd7KsroX
R/mqf+ms0F35juWYE2Ish1mYilENV+dMGbw+dOFpaWSjG0WiE6veaGH2rGZSe91SpK77fYpIr6fz
Tj7PBSlUAL9GrM9wE6TSkg3Mdfqwn75JGENEtbbIo2G7IE7Vrygd+jzfiQG+E/HOveS6BzJAcUup
YtnxHAC52Q72IqIlDS2jssfS2+gSH9uXObZJxSNCXohgu4webCwJpw5KHYKkTqHiYe+oHIyPB/Qu
7V0mkrjLT5mMvVYW812TiUrk6BM2ZZqMFp00D38xIF2vVym+HVOkyYlaf7GASedvNt+33BHjR1ne
sk2pbC5QWRqEPj2Ut06ALTbub7vQVPoG4CaL3/SwQyCjCXDjN89ZvHDBNi6OOlS21WhPKTU7pFdh
vzHoLKxHuY6Y3kSUx0vjJ7qEl63qeTVhSbPEfrgV2XXJnsBITsckGZ7BCWWIxYw0I9TqRs56iRHr
piLAp3nwRtZItU1+3rK0SvWBSZIOuE0cn4Gr6ubhbywvzmBTkSALTvt6OqBp042DQCM0u+V0en4u
qfLE2yv0WHuqlHvHdgX7D4MwruR8vRUGhyPWXjbpzieNZX4RH3j/yWoFpEJSMK/o7+U1WopONcCf
18ZgPytkB6lNiYaqkW2ORvgHO9TNSlBkG0fLi6JVGoOF7e9M1UQ1A4iy3wO8dS3DbyXzYYDbkooK
pWRp9YKR5nHUJQFyu/c8iKOOEQmp69UG6l35DgyHxl7nDG9JqXey1sUjDvLYlUVYUoGPcoM+eO2J
dRANkS1KDPd1qQ+tuucWoVZU2zkBE//khBVhmoKUZ5bD2YU1LaS438tx/4BTYed0q782PWTOIvaP
jodsu78RhVuX6+Iui4mJJWU6eOKfFg1oHClF1+rlkpbngSornJb2VTbGz9VqrKrh01/F6HIbqUXQ
b7nyGOZUw4CbBY6JWUVhggklT0J6EikGcJTroyie/zZ3NE1ozDariH51JBf8xlgPz/YFlfUOCdWO
971jPKYR5IIUJKgi3/KKPeMFWPt/aHXlQNl9vb0lHatPrHVXvIbBMgeIBp3w9FEtZl3Cn6gwSRz5
D7SkYRl9KeVhDNS+3XM8daYHjpuYpx51GCTmWqPoe+/wFS2CtMJzCRciYrhSXoBLCJ9MseGeauy9
LXnymtiOPDET9oYyMRQCXPLvIM1sfWjaOVx7deHuN0ajg7N1QzEPsEx/ls0az5+73FoVCosVbTfq
lqBmA1ktdeKEZnswBpIBmIb2Ky7LleNKKOauoCb51rttWJ3lNow0Ctv3tm9pvJMkAktVCjWopx+2
t0idwnWWxWjUQ+8lMQsOR1wtxle76JuNDl3cF1vm8iwBfuMamQsvGfK+1mbSW8l81qvqoW5p3jFm
Udi/8Kk7XM+86Z5N1fxA8Irxoa0m+02PhAbjWSKGgLFCgDbKzMAOpPLaX6csYO8y9tVjQQe70p07
a9ke9HCGNTqxRcvCWEgB+N4o7C0VILQoHmKm26i2o0Ab5UwqVDw17Z3TVhQuNlkpRsSy7dLxlylm
hemDBwL8aqvTazKSBh4LZqt7VNNwBYHLaSc4i9N3WXd4rHZQcavaw4euuAexb7sRaIfo/T+QBNVT
E0ZdBusG3atElvadKnubHahQfA13wIxx5m2UvmQnLA4GNOvES08zLFMYerGvZ2Puv41UX1zDudBf
o4/SfdUh5Wq2v8gwdNyH/SmGYKckvGPfSpYJ0WR6ih/sY3eN+WRhu/A5RQnJk0BwQP3XIYmxzDSj
5juUWja8kV69p7Egj6kEXi63iHQstm/B+42gPfFdtsSuMCrrKB3/CwnMv8KL0sGnSHwQYxB17Kzj
ZaGf98Gpq1oNTgtmsWFYrHEiH5Of5+OS14GP411KE44/ClpUlybu7I4thjROWeHZASTLBG3AXN+W
gA339bcGVDfZFcNlokJ9t5N2BbbFOhpWhFZiPENbVdMjYl4VQUWV7v4rB/lEiYzx6qMkRSxxaT8q
4Va/oqJXSctY4cfCpjeAUS0+15wfw/TZpCpjFEP0bYR16J1EbEKjOwds7QAaY6sFn2Kk9lbL5XCN
lyGw6yEUmKC2ku0uBW9r9evZDgFS9fsL0887MezVhTWomETnlnJo3UekMjgsG5kEKK6FZST4Uh3P
GGJmQnVmkZQCvwYff27PZF4G4qQVwiHH4LtwKpY4ND0FfW8MFTvavXoOtlG6FCg5CvB4n4fALIGF
nObkFj86gyeyreNYcqZx8XlpVPJLBQ0GvZbfsmeIi2uy1y682tZg63WckzXt+pHqjeieUhEBu6/C
rE+pJ2dSHK8gaBR/dPVDMounvA/Tmm/uqT0j4WbGszRuLa50qlAv3XMA3V86kYrqFdlnJXA6r01Z
j8qVertHVyJ2QF/APg6K5xQTEA/cSIuJto9JqAHEnItXAca++JJ41QvHdF/VzqM22N5QbIjQ7u9k
uAa74oeu94tvnbLW7vnS0smwq47WqrYwRyy4OAiZHYRcyP4AipVL0IUQcP/6Qm9vhYSICwr4FrR3
/Pe6EBp+IY1TuwR+pSzkDL0MLI5BEviceAWE5+apujhY4yyXr317ut2Py/T7Kyg957xGVYZ2l02I
lDhTcNmPUF1IAqNmXHcDn156H5ToTvY4kIsNrE1vN820Gk5inEVTPvSOGFmEbaumUeTHivO+ofgL
dKPDf8XB1J++QLC2RzwLy89NW8sgVRDsQ1a+BfNW9e+G51UimEV30Aw04OdnofkdU3uV14Zv9TMF
FmchPaS2VfKwPoz+d0B9VJsA0Jvd4f1vQTiYNHAxg40g5CGPGKHgArDRLJaiY5niqZXMFflgiLd/
aKxSmbrQGuvMGd4P7rHDo+Lxouklk7cKTHAzJ/Iqhkg2IwwtN59LiMXvRxhhyMeLEOKBiTlX0RX/
U/X5xEbGVmZJiV7pEeATe9m+cgApRTha7vGewjuo0WSZFq+KadTN7dBPHDy1CBOPE0N5Mn28lhAy
T3+L1DSimfWOiXJNY6MdcXsw0z9vtm01ShfFV1QCX4Ebwcn+OqICdSFVqhwydmBkhXWE+AW8tw8/
+0fgNnxLSBIy4pYjl5M1UccnO36WkMaF6Ay25Q0xiSwnegbUX5SCPMhzUJC4kryp4LrMIm1GygGY
ui79Njvu2PaqKLig3M21G6L3p/ss8y9t5FTWSXUMhZDCwVhikklDutuUAAAcJu0nz6xgzjn9PQM9
en3ixz3zn7qWNzScnpuS7Zepvr4tyGRX49eMYASMfH+rut1nwqIuFYYSw7brmacSsxtKiHDax73E
57y2JsPVVOicUmBOyGC4ooA7mj6qwEhBnUo5qsOWMZrKVqiv89UP0AwqVvsxzbT2NAkZb2XOOVcj
lLkYwAHvYEmfWlqiEjUAOrmO9cbb9oqSBKBuezFHGkjzRYIDGNW7sr2ee3I5Cm33z8d4uIeH+7ch
3d+hvxT/A9c6NgFGlK1tRL5PjdlbtbOmBbRU0MXqjix3Lj9PmMwK6aWMuW4qV97qZSogEaZiUI/u
Je4s0pSGJ8W0CY1MLZfvfwS1UpDaDsoMn+X0Qpz2SyuRxdtGh8jy66o4joWGDNf5ENMPcraN2SSF
jA9Ld4SWtlCU0We4+zpEZyzpI/Cibe+YzsNf0DgeWomM7NYjCNYDdU61U1bvoQSY3F0S5x39JASr
fkCyjqtViMjiqm5Xq/5VMdscQ0Mdn9J9s+wAZIN88ATGw4CGOBg25GMejfNcCnvm/dKMHZG1Xm1u
FbUniWCePMmoUjdeEhHmM2oDWqSAcMDHo5ASf67swhCTbb83gAz9qLih7V6f+sdWvfS10fPNInQs
EUfii2c7MdHyzcMgdKq4riXnZw3Q02IGUbi4BRA0p+kstyIELjjoKTzD6W/TLrg9y1YEiHG9lUrR
AL3w4pmPHprv13SAqe1y+KrMruoK23/TExDAaZcVC3NAop4vYcTiU4YF7x5zjQ1lqEcymBtvNQOE
JB8w4J2l6DAwX2ezl/j0jIpBPziqy81Ckq/p5t7YHDCHcAEA2V8jlKe6j67v8UEpko1n4EwSasx2
LPX9GfAYfYkkTYj0wsAV0onRkjFOupzKXPmCFblYU/oI/UhIDmbIQrp+WQZGGs3+q7Xq30qPJ6kU
bmZepV0ylMqhZWaKBzT8UjeoxMnwgk9jfWXNTrWDt6g45u0Jgp6AxbWHsOQFfvG2/7sC+0eKWXi2
V4SproEaHYdrroDQU7zW95rkXMJwwSC1fmhJEsDWa3aEn2rQ4JDBQrjcbDqeDPOL2QgdKV7Gyu6h
3byv7GYpKgsyxEimzCOMuGe3EG3ojEbQZzH48anG0nxQvVZozvbGvP4uKTRdPhD8URnvj+jG55yg
PLeUESad+kUQvz+Uv3SKbho6AnvVwJg2fIULl55ZNRBwUgcKsHmghvHNaedPEJMO+6A2q4emfbt4
8dyrRfJp6eiN4hM39GSBHhXLRfYMgVM11aLPaLbwkxT8l0Kzy4absLCYgSYHQB8gOR6HabSsq1kR
p5FzOLQFUX1Q75aGnx9DrM3Bad2rObjxcmCkTp09dc6VMZqyTZsuCppnkhv5n74GAf/lXgBmKhhQ
kuVbX4cD7fBSiBraWW92GePApC6f1JbYau+O7VYL+iQuEibSlslkdKj9YEbgRHDCu9M14XlG3UHs
StyTf9WChOL9cKADoA+qOpj48FnKwxklpLwbVLhFU2Xc1HG2ukiRaVmGYSodlxLzls0gizyuw0vo
hPxhgJ03qyfd+s+JyUK3mWSjHax9Xrli5GdPQ8REgVTASM4tR8eny8cLDw39by6wpoxn4EtleRXZ
6UeDJ1NHPj/EqbywWcQBJZspVaTCmSJNfyIOjuufNj8o0QDu03zz4fWesfNFZnsz0YFWA6PBV8bu
Odvlv2L1h6pYrwFGcWWrQyRuy3S+Hdp/NpSbmYQeskZ/9bMfLeYkrCZ9dPNKRZ7UwH1yfRu9CAGq
i2CwADuwzGP3t2/IkhVOOMf/bV/JuJI6SPkR3FwExa//KFopCBdPheuR56LtJDr2bdPN9fzgCND8
H77t5AtbZhgH/WEKneO0NEwP0MFEdNcr+P8Km7VEdbuBFY98mv8bDJyRJF29n1G3wmSxQspFh/gL
hz2bnmgP6pV6IN83Yf+S+O2wY45WwxpQXVt0aYR+J9YuhSi0f8gh7vMIUrd8EzxgEt05J7hoH9VU
CPT3mqCtKFZNUufiBuzPxu9aQnqC1Bj08G4ASWCSfzQf6rK8LmbgjjNOWpRXRYN0W6eFfzM49HsM
EtqOJM+3JXFJa5fUIrZrrFibSti7SpkGySfnwwt/Kqea0pAS2brUonuaab4ICi57iSAWu47STnsv
teQe4h3b6d3H7+++hfAWNW6Bd4AuL7cSqfC6nbb3SUJBfe7Yo0dFvXndtA+lFp5L+naaN9RC5Swq
1Nj5/TeLkPFy9430f9yA4pVCr/z/Um2PW29H1T4tXrwKfPAZenvfDqn7CHSqnw/4AueRvfM3N0FI
Sg4jcnxaYrgsXMF6Ro4k0p36uwi4HFLgs3pVjHUtlCfPatZ9Dh9v1CmJT6ylAM7qYNCeATvbi4TY
AwLXY+BrDra8QUurNxdDVSPABSRzUSIeTEZwQJbII9VdLgd18aUMSPqMuhx1LX5vDB/11vKAvDJa
hp4Staxsb5XFbeIda99kZ1cYMsbcSP31DvzF58uCQUCO/iR5SRqqOw05Pc3H1ItYIQy5cwkEmL1W
2mTMvtZQrKg93RkSwl1CELmZCniJqJptJgUNF4J577KLgAP1xL6Bb05i80cLBo2LCe4pvrQosujL
D7WDujbSMt3F/oeQhIiJZeM1ZRe96gnCr/BiLNyH4w7Z3nHkWNBFrpX2d7Q9KXMSRsqKEdvPJ6zU
wEJ4GLqu6zbNN1YFczVF+ig+JlP9jgaXY5/1D/7Zwedtes5nyKc8+3WlYSViDsIw8iHDs9Y8oT29
JJwFdr3kpalGzdmMRzcARW6hFcg+hBhBnfMTcaRhM9uY6gLy+HcxLANYsLZ836UShmmSHeVfBHc7
UW1lXv5PpXwJVwkNrKP42rTN198SUJPsDVtaEZQvIDXHE2/n8oi2whE/MHnyNWcvu4Pjai/2RJjq
ZiIycsgwFkoIp1yz0zFIzkucbzysJSSTq9Vh1EbT2NHq8Xrmo7zZ3+7dbTfU9nTalWkHljrNE53G
07vLvSgH0rZatwcyd9Lw6ACt3qcXO5l8rglNDUFtR6/VlexN/Pc6F49mk8wT22T7Lk78W2TLgzb1
Fzl21D/ZCmw2WILtna6ebt3QKoErGohTmh4zyECu9EnJnsbpSvH2tfktIdjwY5p82eDgdt8zIg9y
aN9PIUOqMK9r1nDyWJR7T+WxLXwF0ov4X2SV6mMpDpCrt7AkB0zvx+jA1IR2VKNjlAIicsl1MdWe
kqykMD8JClO9KLvcvVNJTRG+CijyKpMaTHISQ6wK2jmU5RWRbWPYTCP0yCr/ar5BZt+0cP1dVsyw
WUuqME9UctZUm+cAALrWhLxxg/EO38Kl4Agci2iqAvP+QbA65FSd91PGhr3tM617NVdmqAZZUGDk
Mfd/Q1l89S22nksHYN9dh11f+1sIMhmB0ikXUIyU1QvqZJUfuc/6n5rlYoykAeFo9yhZZuoIrFV1
LhRsq3GD7ux7kb3wmVx5EufnvVtlBUdruUkJO4uvVMe32m5siVsNIZ+TR3sj40KiSKmuWBchZeBk
BYQzxKx6ENKDdafmMOfLTPJVCVCkyikRh+oXmzPgHi1pwgzAUaEcIe4BOyN5b3YSWz1orMEe94Qi
+uRgjyShrH4BH7SaEFfegPRLbEVOftTq+Yeewx0JHJYQfmuQWsG5mmXRetbKM1IpiiXIO/jPWHSO
0bRwMYWUMVT+AmBGzI7TI/cLKFKoLugNxtEB19wR8EiT6u1/yMIuHjsQ77JuE5pXWmyS8ZQAAmJM
HN/a/UpT+uJD9D3HCXDDmIgcN4xWKLVfCLPFY3kdHoAt+9UfLVcodrdVfdNe/ntM2+pgbfnvsD6B
kH059hSU8iNhkT/4ppE0VO+AhEwvQTBzOPuZesd2mLX2Lp/25maWs1lys/Hf4uSmTHIeK+WthcGL
nJQ2ZTnV3aFtCsYhsERZRLALS9PMACPLvKpFowbNcC95B8WV8KysjZIhwxzoqKjiljyc1KdftSG5
Wfv66dpRdmiVzTrzkodssTXTv5+8bEvNuChaVk4LaW52B2QSTJb9gNHHYPQLDIidL9rdpdFacMRT
AuxGEtbvogOIoHmNFq79p2fMF9Z0xO/uuyBeOofdSSK23gmxNi6nJlZkqtlDSDNxI6AycUaao6NB
lyRI7mA320NXtc+TXa3XIOQht4qgMSqvAgFe3DkjOCgH19JDsjQEqRXc1HJ/lkWy9MkxKiVP0nr/
KMq9Gie5vW3l6fgRfLrauJQrP/EtP5bSF4McsyW2qLI0uSYpzZCJmD1tDQc8MNrGeF9vKSPtOgge
LvTNZTUG67POHnqvq7u23j8UnLss2E3eZpOQAC22om/yOs7hj+RptOl6MOeW1pwMJbNKDTCaeFQQ
dzd+EStdbQxeMYeHf2oVtKSxfhFkXP97hie/x9MITeCFyjLzM1a46jc1TfSxQFC6Px8BD2jh9ekl
S280FQlq463icPWLcZv6b4R3GF7TZ8wUENsejLofsERUibEReEOCwfTfcB9bBhDKLDI0lQD276aa
x8Y4ythP2C9HAuCh00E7DZdI3iP9P+ea89KXCsajp5h+Gg1WBMFMjICXa1U/wXGNkm5YScw1f2Qw
o4gM11vyIwSQNqv7JCo8AqqbFANx4eltMC8h2EBM+C96c+HNRTXjEbT9/6xsCO55sIZSKoB1RHXs
IN93rXeR8+3oheEH3OP9KFZFqN6vQpgMcTtihqZ5VcC6yCop0Ud+lq0SOMTFCL7QepBj7KSAXaYN
yuO217WHi1q8bfLEiCHCC6LtfMpOw8YHd1LR2AFlCif63oKaL6nIJp59vEicVW4704Rwfu7Jhl7a
uoAnkB/JWW3wdxTwc8fD2lrl0CjDMOMwQU2xD5pE0LmsB0aEgoYGoPxwfxc1tQYDJVJMADMUmhYZ
t+UkyKYKZLjr1WD6Iw4mh7Zv88cZ9lG1/qFCcWbAkN9wdxpHj7+YKCdVtCZ2slXYjZYqVSlQXO7H
nYaNAdTTrDY3zJ7ubjZ9kJeMRkkthLIXBGm5h1+ta2XlH1fu/dAg/MWGyp33a7DCicTnt15sDpCO
lcUrUZdUTpukB2b8wRGYrRWAN+AgisAQZlWZI/9s/74H5w1dgAB9BaK6AFmQDh0M/RsQQ/9BFe8v
y9/EIEgpXh9W7R7dz9VI7PvPUmXfHteqTR/SFtf1Y+/HhAadUghaNG/iLU8IcSNFIcjVWr48xeG/
5r7XAUTsHSNV278j1llSFCIyq5sY9ZA0JiyLHPOOLBFp2AMHnvEnVlJEUqLNQEWX0NdZ2iS2tSej
widZL+xD2o/+6dTOk3v/qVkEr6sRqEjJD9P+FJAzNuYVddg2HA3JL0No4rb13GtAUldEJ8jkYNnl
Pd1GF2bKoPHpkjlxad8xES1MwuEPtCTHEkMqbFMg6bJePYMTd67Gy0NyxMgJl2PeIe7LcLgMfoyu
sKGon9KFEYgjOQ679f1CFMfvee7j+VSYs0I1038jsJ0npoKY05e4oe+kn8vdtczD1okeXbDA4/pP
jDhn/Nt369l/Exm/JWdmSQG5pfW8KVwQmhr+Cl2WBC48Sby2o2bE2Emt8U88CT7LYklXBpvRAdH6
BKvWRbSRF7YFPPkgVF7spip8wXU9hlaYfTRFbrXht8siQF1e1rmj7jz8SkPKoZEwS1QpILetqQ26
DD/ld8IxLGEXpYbATsRa0P1gF5684PP7PIgQ6EhMsKm5Z5DfSqx4I5bUQO2vpGq2J3rhBUrG5e3U
2voKrLurzlNMgE/kfPIFSLVjBZd9ansPmYh6oBYvXif/3dn1BQljkHHwGsbpegTbg1TgQzru6yoZ
mrQcAmdwVxRQkzvgx1NYorrqC+bXe9/vw0FvI3+U/YXpRvPikhMPG40aPV7sbuGybsQEz2G5aoEZ
rlyWWvotNRBR1B1VpMm989uKFHByXGBFIUM8OeT5QHoDLHZeQo0ZNfdk+pK5WjZjSVv5dEYTKTI6
0F0zySJJHv9o3hgRX4d1XVUqWoPBjvpyOrB7eH89VhXzWeKoVdVaxcUfRZhSn03eIMSlt1CgE/oF
1s+KL52Dq98i6i/qYLW5ISKHw5v/gFNKgFOQTiXzJswAR32NRgjF+2mIJeK5WnHa1LG795loDjBM
es+G5qscqikVTM9U0TtzU2BTifCHnlpPijW43skB3HTx4JkRe3BYr2Sp57iMhC/PHC0+sCjwx/ik
4pEQxY0S2K/FiOeKtjsT48kLig2CyiKv4KO8/0272LABTAnghYMKwtDmtHhouBg56I/QKN/PlY2k
WvisjAOa3cREsLHe9XKP4HwqpIpx9rd/Xs/1P+d+n5e0a5LHaPqtIlB/GMCiJPGu/CRr5XxxJMX5
+dI2Y+TZbDjMcLAuj2J0RvAQqiN+DCYBP5EnJ5Cuvma32mQ6ykRYM0foTBxxrzALkW7mB80We6bq
pHvGCGf/wagQJtbt9ro2/7+86Yjo96TATtlvTTLfENsWTPJpvkV0uB6xSQOms1+CGUYx6fCT9OTx
PE/Aw3ssjGt18JKEl5zyWUz3Iq1XAqvKhy3WZDTxax+nmiFIdWqZDBaZkf1BrwYCe/yqxEOTDDww
WjWFZcD4H9ld3USel63HK8jf3jUsorDdKZCpc7IhfNAXxZMqRTPwLOekS/Jv3jNTwCIMWJpGwwVj
Tsg9toKnDayKFlVQa012gKWf7nGN+u0skcBRY9kpYkiGUW+7X67oO7paN16JQ9MPWRI/LAqjlcSE
7xkcBwznTlpPODoODCxoojzzMMsoVsUH3GYdAdsboM5acYXPMOprf8lcMWnrFIEbD13LGtvfeUyi
BvaiehOXU6ugIN03iQDOwrqzH+JwWNBhkKAta3OZnm97mnEnRgd8+qvfUR+IzawcAMvLMQQi74AB
+63X46zlIf0gOPUuqU+a4SPBdfd+as/65Gm1Q5izBxF3P2VVM0/mwgM1q4zdpZqLW36aq7iJ8j/6
+4EAZO1a9TXnKTsS2Kmu3ve8926bBCEUTwAg2ty3M7TeoOSCsx1vHgc9Oc1317h2q3/tWojnus0U
YbzYeU6DiRI8Y3CxmOFSG5VfdP4hCj1kwempr8tsQwemSv1ksM6CfpTT/cQN6dZXkGix+66MJS2u
IF8IpsCzjj9GxM/V/qGE5CCgEtQbsoiJNS6hVdy6vOAkpTDxja3ny7JwGO6dFquuH/33PxuKPfhi
4anxPzQztYGjcGlSIQoDrGXdebpDL29Jr4pqHsR8WgJ1isPJIPytbNFO5ZaxOKqgkErbfcoMtso3
kkcpe81a5o2ReWgnFK1gQMnr7bwccqvstzMt9+ZjNrRnYgVyyMNB+yRa8co4sKTr9K5H33r3vE0A
fgQ2OMK2x1QnHSHxqdZRaENSIuVxQ0fy60lKTt/B5tHlyOjG+HPv/lf8zVQUoFyvCk3ytgMAvJIh
UIay6InhqcT1lYnz47f/3bXX4wz3hua4pL9SVekCF/kzO7TD3/mN8g+S22uo1KyI94TvEVfzKIyc
pF8TMFxgI0fAYmIvWr2pbUExH2x+mmvhq+L4nNKzEqqr44GrrgfhibDDkYctuVWeLGRuq2lSwJUo
JqXaTj/31DiWR8vtFg6Sy7D65gHLRqYFddKS3l981uqrv5022SXH19xcfp9wLxw9SvHzdeV/Z9PR
2sqrbNwQj0LFYbVsI7XKO8Z/Kg2UcL3y/6LfRPVUudixgeT3S0XBvvG35XY2RlonOScxPkLx86NU
4j3A9wxSPGwuqs9SJlrGfJbHON5fGtIvnbZIjexCfxlQkUHOYn2XUqg3OAf0JWFI3S1reg4LJmjX
aE22ESspaqgjt3RtN7DmBUDBzMPkE2XfPKOftZb++Y8KDvdZpEJvgrzu3G8XUPKCdavoL6bjXfWR
/trtIcYkl5zT99T4lecxxXx/wsOqN/UWQyFyTRRV1KzgPAYyZPNe9ohDYnh1rySWXVDDPNijf8ek
RC0832rPwmFN4h8tXoWpOkEJpoSJ4Pv+tH/JkSyAn4fm3t1hpC2QWtwEgPF4RGmzjLiFMzXaX603
1dW69T/yoF5d8HwpU22+dJ1x9orVDI7jvlvwb3eVmPv1zTwFe6HLRQrHyEaIT01xklyNc75Wmw/q
JedOf3jGX5cR0aINjOR5lOqrulP4jA/Gg6ncIdAsmVoWlVwG8UZog7tIK8hvp00O+Hh8O94YWWm8
09I/AxtEhwIdkxt8dCmsSZi8LQqWorXk1LYHg0Ba74Zj1zQjKt3TjPMheQn9GMxkSm34DdfJPi62
eC75Yu+tDkraTlJgJw4KyG4q7nHyctRj8LFZQYZjylruzBS/o2QQgTizfiDmfc3vUbyhrk3QoZ5B
eBIxti5IKeqMhbaNcpOpcKYtIz1pw/zcWuKAeCM9bX23gwbZ1Lwt9NmRyb+0GO1WGiP3nQP0Fa+B
Nj5X4uxNAOikDz+ne5svPiSiHlcleOki9D9Zo8K5BzoNRzyRgkV67cTB+12U3b0aNKuT+xd0hX9Q
qYqQ/xtW2ul2bh+OWbSNkSiDazBRnOt22WP+1/06s7ggJxjaTeW3RwGMt6yvJf3YC2vSynoTcQH9
DPrLqQ3jVR5SLi2c/NNZ5qQRfHe3OTpFFOVGnUl5yj6JCOol+bQ6GMNBBVFQVw6Uwzswx9q6ZVlr
JHaGIVo1EnbTqi12o7jS3iKAnQTTepvZjEdKqywzfu619J452HQYhjsZH0mGi24fTV4UNeuAIWOr
Yfz8fJrfQywL5SoTHJzYifyrYu6giesZBUKGDcLGejdrfdlMWrSrbuSFCbFelnTVvZZLXpL95WEb
F9TSVXY906XzaxYeRhHvvrT67xYJHCgrXaD0JleHvTwpKPdLko0KMNIxzCtTITEY9aRsCZ0kSRdm
0EB02J97AzjoyiZkluveXqdccdgiSIDof80t6VeZ7DR6P/nYBT6EUEKHF3dwdWVcXlXzMpsG4Jai
Q4j0JJHLTNiZatqh4w6DYsFAi30hDV+iUPvgy+MpxD9agPVIcGHfyI3e+mdqQzh3efESWq90tcM7
WxUp06u7jn2P3zM1IYpcTkBXINzxbDJOY8Qgborx2AlxNwodWlBXxNbyv5caoG/sCVgJUDgOO29b
QefzVfvFuCkxP6vbn7mEfJSxfesNfLT+5bleiKPDbA1sjN+aLhE0s8BAKTRrvE6P1oL6ANLoLNFy
0oIDvWFrYzcTca55PnecAteN9TdGCxe4oJYJZLSR4o5rK0JQt/Sf0wduRcJ/fEWFRGAlspGwVtOz
8p+yndk20XcusFfEP+dGQIWoIUd2p/pWklAfOL4Yx1WZ1KvUUzw94fmb0Ui2HMVF5ZOxaqKC2fdA
JZ8dd//B8RKOcpqtGlXRyvCW49KiKAm08wl+gD5IKVvpTbvyySHBQ1gW9A6R97T9Yxx+WJHtrao1
M2IZdwtCGDENV1brLrykCJFK8ZasUxV4Rtc3qnvV/EMfk5A6kUN+FGAjHXt0VMfZc3UfHOfsHdj3
M7SdH6yDE+UvC+ER81vzVNRP4QJdweZ2EJKgSO2VP13lGvXQ2ZZgiDFZSLyDnz6xdxkOFIrFvFUE
zml89CP76+phnqM7C8X9McuzuwFN4wVj9adIShBn2d0hBUHeT/UUWmXou7r+QE/PrTzwYnS6ZvLf
lklG2yf3R+g9XNxiVXAeiZmV4KNNb4uo6UH2DU9PD2I/JyMLikvZ40Fyry1GwD9JVfKgLrlHoMkq
S9UR/8XM3+BWGTYWUNhNAqtdcL3dsgYUTDST0NDQLlgi7WuCAU2DiDwZF2Y1WmT7DYld7oVNk7ne
Uw3EVjusF2ZibwEuVL82oiZ2F3obQ0Y4Hfa3efKZa+a6G5n9o7/ex5GQUjcPEI1yyhkrGseKgM5w
ucLBBOJNQjrSXERv55tcfeiO+EtoZwuV/KbE75s1TMWDa9P2JPBPhRcISmdgZNi33ghK9/NlGaN3
3DXAH8ZDWGAvPTPvqFIRmth0PcN+a2s5QsFC90I7kbjOBU1CyGuagy88WSaIXNwWIwbdz+jxAPOB
AdRPO53ujHlM7ROjkxdB2d6DYuNroP7Y9nQ+cQWeeS0D/tmJ9Z3VPeSSWT1XJd0Ysm+5jMwVUozo
Ox/jMps4NdHNyp81eDuzDhjskJOdZET5P24NPFP0Et86gIoUkROOT6o4OB5VhhQwZ7sH6pGskmkf
4g4okxqxIy1eBCkWJ/XIEjZEBn0NPCVLOIubD9FhdyTg/JsIA472bwSk4zQNQFvB3Nv6UyfRrM/l
4fGlTctLnQ3XfHdxNdmZIx5YVxsA40PzlUMO5Z3YchIjxSnvY7Hn8yzr9ro/X8VeWr84ZW1P+Ceq
WBioXPD+0mEqutNzedow3RWpGXFy7EIFT+IhMzVGDVI/Kc69ecdE1+XLnoLxW/LOtOaHK0fedpFS
C2WVv0jmcDZ4U4PAABfSsne5thfBaGRNyGX1Yvbkg+jdqybanGX4+Uj1f1PEZjwabgCaFzG7+GhJ
2nteti5hfdFVho/7aZs/bKT6zMNqSz2/1+lXwYts85/ffpMtsyDBJjtyqU4yNfW6+kcseskiWOhe
BvRra3a8dsVWhXN8PnHUVWGFntN9Uytnzi2iULzIyyorY6yBU/wU6VkF0Ua1t9LK15RyqNSTXeqE
HYgLnAG60l626B/JIRpeInFnFcE3dB24A1p8gz2vIxn2cc/2HBIN+bcS8rglAnizldVBqbHYbDZe
ON39mW3KASRO2csS0tv55VjclzvvKRvzfRoFatJPotOjnIBZONr9KKdyHfxdK3wuusFApfYwX/qh
GHeVGznb388EzkWn9+pcjPDQkj2uOK6YQmsCJx8K5MFl1aMXJV30iU1au8IgCCIhC4AOlc0vOXEV
27jU8ApRZRUewaGdTOnrkQo1wHuZlvU8ZWW8oOTt5VDyQXZY+XcQWyZJfdY1GhXnn2BJhucOZ5+j
Mk/sUroCHYYnPObYaVwvyi0a10LdhTAHGHSh7FmbrjogY6L0nzY7BcVzk57k+ntmyGOdv3Avt+qN
ghhInfgSEndruDgoxC4K/S26Kb61kqaGaCE318GAtjF5baJPj7vWfTT9FZPqemBQvWATPDtNtaLG
ynF4sM0J6MkMQ2KNk1TOj8rzLH8AaBkKjFaSw2MUTuO8EXWQLOfedfv19stThkPDmihlZHAf8GSH
2RxCo6gfA4331GIcLym3sXcpldp3/gw/gM1zl6zTCqAdL9Myp12J+irVOHcfM2hT4E4z/bSKnEZa
JOwKxbfeG86x4foAVntJGJcWJEKVbY5rvaxuDma8BQKsCODeUMRwjT0Rg2xF0Pvx+zZlKxN+3n4T
sRokkCPFuLPHVGTHHMq+eet21OT4DQEIRm3AOQO++oHp1IRCgKt0ETiN4bMLaHVO4HmNLXAQaNzd
TdbOSDYsJM7+OwArkYdpz+BVvXxSnZM8gJQrx4zNaPu2tPybudO772sLgyAGA+J7f78BH6KaGyYd
+N3WxARfPJ7pfR9tLGWseWvryQsxmkE/Zq+bK8TDrbfzMXkAgZKngqRXNbtp6zTHt5JUdg6W+0pF
TDpQ7s5g+2alxSSfwVFXkWbZSdJqEeD07g7siwaL/uEiMllBCpPNP6dy6XaZ+0ggxvw2U2wxC3S0
kLI6VqqUVt4HWlvALy02Ed1emGK1z+gNzOhe3rX0SNPDIsOcHwmQUG/fr6k8MHD/GVJYi26uimio
DkkfPHDSA7MJ5mP6DBhdb1LrDo71LhJzZCxI0wOF5ADMTibjKa8rpZMzKZKD0/QmOf0iC05BZauk
hAnPeR1wvfP5WbMGMkzOXPhV9P8U8L4jpiWZoQblqCaLfA+j4ODuZP7ezlpxL9yBctCbWXYHZCkl
daBOWV5ZVN2VYNRqqVxbW+z30G2+z7ywZJebFeTjGY/kmfUkOjxz9EM4dRXR/2Mk7pOSscFswS6W
S94UHfI4z1YqR8t/PfPcXN1R/a7ectRdS24pljNG/eRWUWuMthdRfOa75cRGyTbwKQOCvCci8oqk
uiqSOqPnOGunIab8+9ePXKje1xcAfG3LXsxwfHfF9e/L67oJ8tOaf1q57eJ8QBlbeewVnXk6hmis
qZ41qV9wucAwMeI05wbgFNkhuTz6mXLSZqUixOULPodt+b3wqyeV1fyKNcdqoTTtEli4/UQJc7nN
mbpnDtP65ngpTSQNq0nIB3PYFxlHIb3qdGuf2P8zY0ZGWdHVa7SqxvBom9/4P1K+hDZDXbruO+97
W+0p8aBgbpi6c5Pa3267c8qg6VEWJzsDJlCc+X3btmXbTjO2ed+rXx0IZ2ZvpsEIPd0g2GzcfYaM
zSffuqpiKgfzTzY7fquVZPhSjlm4BbVMPb70CT2SjneisN/VZr+LlPlbD/SCBbuO0tsK+0vexngj
lIU6BC3lck1vKa7zpR6L0WgIRRMkm5V4MGc5Qxaeg4ehMemWfkj7FejjIelbH3k0OIbGamWfUode
Um9r2dNx/Yjt1+a3GT7t9EuChAG0O5jXR+AH92CK6FfcLDOoJnMZ+lUfVWZYr3sr6Y/dgdE4i9g7
KCLrAgtcvnkgV0e5h4eHlm8B5utcbfqfFyZeOCE3n1D4MkBADLr1DIzH1J0OMS5hAUdUq5I7S6pY
Gkw4dPnAKvUetQTTXukwApyNx9cmh7U8pXjasb2EO8gkHX3o2hXtyv17qB3LkSTFUr9VlfDzG5qQ
nN6+4Gp03nZJSZsiA4MfaACv7pdcSVO9uW2HjL/ERN+T8HxYvFJSBIz1yJRciua6dH8c10v7ewAp
86ObxzM5zjH/bp5zmZqmvIAFWAy4SvzCqsX91IIWsDiMG4PQNX11E09BXm77GvxjrMsqGIMxtxrC
W+tXLQDGXIp7NsaAmqgPwUrOFl8/A5G0vgB0z6RieYupWzYvxpVr7yGnEheb9zxnO57txbWby04f
U43EP3qtoXKTcXR3n4pId/66BpJYYbiioVwhHrwba3Pu3LhzSQopMgTWKUmAdvrQYHopxy9WJ++V
pUJ2rXJdIe2ncJVQt0RDjgd6v3ZNRG26qP4y+q1rlr2/A6OsxicmZDurrhUoVsNpF1FpbDGUS6Vq
3DHJ7rexylabPFz22j4y3Dtr+Oza6jBjpi4nyOZb1ZMnW5NawtC1mcgX/B21vVNtt6m2l/VJz2y7
kM/+v+gmjkhuozODJ/C3sTTm0EhAMI1+ErGILBa2nfzyJfRrzPx1ObQY0OwWSwP4aOntTydh/yHN
qdd0fPNMdcLrPZFRogxaPw/4pwMDnkPsUcOfvGgg6BoCLHgekcsk+qLZHwVSzBOfLOfJpTxshI05
pJ1rRyu7mbomQ3WQsqMDM88hECjvE9ZOAeQEeXvnyhEsy8m45H0mtbAmCCjKR/esAt3gMMloozhD
OO9JS7ulKUHYY0e+cIwlKXD1rkkNjtkE3gNjjYXBqTnbj02+ijwfSV+ee+a9nwKq068DVnTYhLjJ
atPAS0lqz3PRW7Z/evPvzHsBsDG9icnYmMKAREoKBY/+A3MKbjnr9d7J6Dv9hW7cPFLqX7Avh6Sn
pQ4rLcoMva977r8/lGK+nhffESes7x9WF3XHTgmjz1XIIQeuul1RrRHuhj5u/tsEoYUHXrKaD7uk
k6isLyKUPLHCZSziqwRjC/KmRhZKsz2/pFy8508uGG5Czp70jm0ol26pl1rEI0n5MMp7pkS0kjsu
4Dzb1w+qvF2T75J0F0624KdwXmfy2XUZwcECc+BKnRNENNrm/b1yQ2QKdhwVaJF5gVqiX0+Ojg17
mo3OLY9P3R5+9wLE0YOt41k0zNqd8ULWZ2HUsHg0VQDfswDgUlJm+u2NnJyBmZ4N4MpdSS+t2MnE
W/8OqmMS4GgWFtUgvbomJfTtmTA/IhIyKL7NdxYfVBgkWsfoQ9X0blZXF4CaBaTMyEmP9DPviKAS
APzidbxe0DJkRMA+n1/f5zwi1SywYWNwx7GvTh/ohNGC+S8tFTA1vKAqcIQI0J00+6E6CB5z7EzC
D62unIUEM3lsdQFV2E/AHTaWkhX0SwfZJFk7NYUNKf4l+dyoOFBOaa+KO2Jhnm2No0MVzAjJsEly
IcCcMB9GmwmWUU1lqdC9k/9XLCmrmc+cjFLPDhQWnFQ+C1ma0Gx09kviTKw5WnKSaGqo8fCxwOeQ
NAMmAtQ+d72HuDIDDcztgPvEIUbMXSY3uXJ9MDRJXM6M9Zz3KIhQG7TQlvYacjZHA/r/HCqX4C06
vVDCDeF8t2wKWIH4dJqeQs7puHc++Rt50NdsTMptvjwv0UE8dlyJEhba6SeNKI775O53b6ByEDm/
tRTYPubFJHUJTLJQIVfAcB4MO305Z1+390Ybh7XhpGyEThHORVi0ue71HjyzB7ZRilKIQ6SWb0VA
RadVVbgxRm4nzaAHWRW2dlXCI+ikoWdPVfP0hNCcwzBrSt9seGK0g0Fty/zYIqmH+vkOKqLJkrI1
q+/FH8YWxf62D0uTn96px9onA2HbJy1LtTaty+XrW/jj8KVBrIuGGizGOIvw0cMurDgNAuwprPP7
c8nBZ3DQuUMbGrTzgmhSvUdniid8nkTlsdVBBJhjCJUmaBKqzx8F6Jm7E8QqVQQ83TqZbD3UTi2f
s6zr0rsm29e0oIpY2gjijd9odtj/kqo5mpYWff7kq41jZNRtvgLYEI+9qj84C7GwIjQO/5bfjQbS
3eQnRp5r6mjjG+p1nzj6io8T76xIfM3Vm8TURVfovmhq1JjIl+P1UpkO5GCK4C1OCwJIwM/uO6u2
8R4fEAQTL3IUPLCQs3MYLREpQer/IzFlkKFhKsxMCa/zNaVGhd2YIDeNzN7Teepsf+oiJoFDa0E2
nKdrzYxGrQEkTY2HRjj3ZpZik/WWKcwhzC0g2UWCs7FOlj9gYLDIawI1JFhWrqBsg5DknYH4Bdlx
JGuSZ2xcJKeWnv7kBxyqvojATBN4/QPmR2GScpLuX58o/ZW3On39pMZcXor2Ux5gR4KFM2UUsfM+
aVXeMdlZN14JCu5taJyS4GIC0DJ3w6DqT+myMIce2WKLEw0uSLL2wbs/QLosY6vatCCbVKHh7LTR
6Pfu/LANvwtIEY7cuZAOvl0FMKpJc6DWl3/yQzKDf6ER9+qe1NKhEK/kJideXfcvy+aJB7x5PWuP
yWJHvAcXLOD+B3s+hs2nCvsbUDGgIu9XMakjCzBJ1TUTnyHlkvpJ6vmnUQypeC640n2dVFGkCbO1
p8TwRtARPG7ADzTcqzXSXZx3Sxt3tP10b037AU0SO0rcQkGA5trYOAgSOjHDKOjJb4T6C5ZpFP1M
LkCAmWedFRXqG7F/oHWs2DldWjVvujcQ/V3MEP3QQYrkWo6FZXYnJSzZ0x2mmDOp7rj/FkUCVCIn
QWNYczNuGCKREEXZRzodl3aTdBYAhcjb2LeuzBHGbojIYmkEcpk0uh2y+2v9nM0+QkYs9qQTK/7C
rky9ghTwggZs7/lT9HoXH3rl+Ial71gSPR+f0xeC7up4E5YA5EehTGg576M78wdpqFM/vUYTpHej
4R8qUZd1erkPtzimGqtwoBV+zwPX0a5zINhVg3BlMZWrjFDm8eUEjxo6/p7ENoZlOxz73PEV+jv5
Tyq5r30LsO+624h5l223yHOVCk3QW1NfJWEwXYFYitMEFSWTWtSpeHWHzUplyYEeYvB5WU5wB3Mx
jtAIwXbT7zSm9cNGwVLRc3/AFnVQY4g2ApT7Br8XevD6T90lKmGPuu8x418Ur9bsvWZtNZMRLSKM
iF9OEi1qnlEwM7Dr7WhjXc9e8DqR2S0bBuRF1MJXZHq0jzbGfL1PAzQJXRCpEdJ3h20kIqiVWk9q
xTUK8FXL7xMT+RqLk4w3VAbcpfZ6Sb/vbRwhYyQ878DFkZhF/7EFCr7TtZDJrEeSVP7BNtskwZbR
yJT98zBT7ygr3D3+5P39senkq3m4gaPh6sK1IOTU6JAejFlRAivz28g7L4XO2qJUKASq2QbfcVQg
fpvfLsUQzer9rLlo6asPM3fO6l+4tzMWXYkdR7nm5j/GULdMWp2se+iWi2Jn0w+/W/5htDj0hgN/
0B2NCgCe4QIh0UtQa7ALF3lfRE7acy33nBZBm8829SQbuSyDp18ZPdNB3KhegCqP96kg1d7h9Y3C
aOCL84LxUrFetAldfWOCNTqb5Y7UA1lX5KK9HFOGoKHQkMTOyLGXJK6jlQpQSJHISuC71nw7GaBO
Biw/ijJrIsak33dBTAqzNJS6EacvYTy1xf/kX69f+6u4WmZPfLKOwz8Ljec4053p3s3noDXwXYPW
Cxq9yw+6lRY+Xw4vpJEG/PZzlgP1TzaB/1dalQt0lnv+3JiiI+OTuNQVWD70l7DAtLTxAZb5w+6A
7RsWZO629rI03/r4QmWIF5i0XDN8NQSnN4k9YK2gipumuy9w/+NPvP0gSq88FVBmJjmLJr0s2a5w
UywUFGtbXg3CH3R/3NS+eIMCg3/jfG/hE1KK+fNv6GY8w129jUy3GpIzVxKWbv7RXUDc5K1ilLIi
Q20clwtxfuPbTQ9PK2+mFe0ihdXojTKK8reGZCxJiGLlQhHr0BuRb5zTGwafQpb7zlgapET4X1Fo
QM32p4xnwGjiGi1yoMZzZDI8pyjAdlGmAOOlaNNTKb9XqNqx7fl8n4/kTiYwLm/0wbOJJvgHx3Wj
gqSG2LVI9QV/jW3AEZypaMpPJNFkvs/8OKeoEgnMakv633ZrSDK7Lhm28pnSxOCNrHt4TnFYeqQv
ihVkwYqeFbVRbYrpHwWmsVrPbueFvOt+zOMe5yl26S2bvj+tvUvu4XAkMq4OgtzfOiHlUe17ABXe
hFS9fJpb5LWBYadIFp1ULirGNHmI8ZscFIueOPk1HRJucBYh0Bkxq2OIkK9bsUpvsGVktyeh4ZZF
OXSl1X5NdCUGO4hgP+NDwHDf8j4tBMiJAHVeFLSzt0j4PaY6WbPoLAkXPLVp1Qclw9uSEkd4AWR4
dwBIAW3uXJN/b/KFVvR4tLcG3uRG5ql0x49DXoAARMGcNYNu+v1hrMrcBZnDW/DPdpeTQ7BnIqxA
qURvjK+XCrJnEgJOMz3rWMpJWcaastXoM5zAQ9fFN4lXFX3HkSspCURiULJEN6ZhahQQo1Mi/dIN
/c8cc9uSN+kNpFxuGbRQAG0o+dSns/VQutxOGkfJy0uWVfssKXVMbe+SW274DpQGftKbLq2MOcLa
DeFHFAxPoYll2j263XW3fujupYTyxMXEmoHpiQRly/aHi81pVksWjzwHW95Ah0VAAxkHlNjmMcdc
7qsVfXFdkGLiikZB832ieWiiI5IKznjQPpHPrV8ooyGOnxQig1toC8FamgylX7zRW/RILtkiUKVx
fVjfWNOk7kaJiX/LKDuX30zHJOSrdSnoK5rZyUrJ48i8zW4aVsKujNi+nLVphXC1IfYDoPPtcsla
okb/oUE31vgizgHhpRwemY9VjEaik/M2xjoFZAWDs2Y27BpJb0VQa9scWNvULszUdxpd42dhaZTV
mYybC25Wjrw7zuFJkSYUVKMNOfbOc4a3VdDgPi6k+m8/Tux976zCxy/7hZs1vfcxMqL4798Uk+gK
itPuextSGId20sYP28TVeYx4Lze3H9r12Z3M7ACJeAXsRF5iwE+cMc1AjKgxpbdQZiIpzi8JdL8B
ohq7UKF8q8xZAME8QdjIRmnvhYEVBceA//QLsnft7IJj7HeC50YwtKamkz0MV4ltTR3289hOizRJ
S3K3jV0HmK14d0WQC+SWsp9lXrl1RNUCQ9UIYpj6uhqaKmsbRW7/CLYlkOYbCmkvL5HHKr+5KgGx
QOv5B9TzPxFmwoHXhEz+VsmRh/3ZAqUFhCV6odw1MhM4EDSIjr2sdzrWrBELK6rEpLMSB9NiBEN9
+4fNaxv6TE8WmbG0KLZ8KYPmF8iuVKFCvblDTlT5n7iALPuY5tjeCcfJMktqhwZQjJxEVC98x9DI
vw5uuu8QH8F343LD0Jt04GbeIo6vQVQ3oqfLd8uYoTqLe7/jwWjq19alDX00g2Q5ZcK/7iKL97Ra
RQzNsPeEJfD+9chssg8JMiHwTFGxCE3ljKB+hSdpnpeZ3rP9/ERz8ZPe/4Cpnz2B0R8FKtZuKfFg
XJuQlPt5imP2ta4kfFFucxxZcCmcegWm2otTfisR58nD4A+ZLJvcwCVcXBAcniN1AHgkzz3BJmr9
aumTou36IJ6SE4caDgPfpjYGhTBK6Wky3CgjVWfxJWwSkKsmZcaC06ZjVnNgfEmNM9O2v8xDali8
xbLWMBO0ss3mYlh/rkGtAahtn+qZM/TfBVebXmoVSehhWYmkPDZqp94f14qnxmepuClOgdi7pQd6
HZvrzCnq4Ds2ULTLNVYzrHfaekESxI9viHlM7Rm5c6nxv/RL88zTDOJ5Hokt6dxtZAwHRqH9qJHN
ag/lR1kdtb+Z+Fm2S8rp9Dkx91yMokUQdbpNcv3FnkwuEezT4cRYIEqnDvJgFyeLtY+9MEQkE2FD
0F0g2LYgA6aSd7VfLxt26amR4iMB/1+g9ZByGFnqOcIsMOnmY+VyEc9MtHhaKa3oNIhgi/5CYMBA
ByvhthCqioFIZTqEJz/HhfVp0cnAQ/rjV4++2RaHL1+9ASbnhUgtJkOlZSe3Mlhc08g+lZWiMSs4
GG1WvnXSIXOQ49iopP35LIkRuNWpySCsB4NW3oajtfDgIx33XZP7LenaIrAxNBoLTb0slX6Acynr
1ETrlXDGFIi+U+VbQrE6bZq6J5cpDEWepW1s6kHvzK5oL+D85m7cZaGSpOdBZ87IGy68V1qcC0aV
3HONk5pykXil/xjbTJOHvZDCShFew74BRBAGZ5oaRrnV3VooMb9VVgfT1c6btWmdbOzv12jRTqGv
1renAbX+TpWmIEgsGjmN6lwI9lTf8CNeztCrQpJTPClQzz8x+9lqzqFcZBgmq/z+y7DwZvFf+xzX
J0h44kB1G2EMxJy9wxUDu3GQSYwVg2ML70v6bph7fiIw2LgN8unBvOGWYBcVPezx6OZLxLJMCiMi
iVMXFmsJafxuQh6tXmlhVK2jNn+V9QINRBtsAUqcsQL+oBDG8UcTnbp7LqfWLE5oSXIb6UBbjH59
Q2GLOd1qEw4xyDbPuaTCriH/buTU3hbKwUz+kereCOErcQFjmT3u2GEmasKBHoLgrDMMjfzh/qkA
pdJ1iuwC2sySothufFX0x3twCEjZkU7dCM3JF/PUsIf4APBevpVnepmkySLFaH2/jpOl4swHsSIn
FfN4f2nTH6uHxogkoc1YvLIfnZRZod8MvNMTiwBuvnrspmG21MhrWCf1DysfYFamUOStU6OiV9dD
SDA74ORYG14pJ+nfDIGl4mwGOvyw1p8rBowiBBf6N/sntdPGyz0RyxP+/82mTF6G+uXkiWMKftQu
KQp2nE6zE36pcEkMGb3xLZ5OQIT+xkafAZccY8e46iBdqlO+iqw/omrDnON5N2McL8o3JiZErqqL
VDeLHMFV/0WA6bMr7QW/bi/lxMh3gAY0DrIv9TOx03DYNEdDUZ/rPVg+7D+8qsKef/mF4W3oQ6Fk
Otq1SNFLP6uQTliVmFV+smBIqSuhYy20lHSpq2vY/sZfcOSDXDXagi/LcoPos6a/PNcNM87nzIW0
YBYNAq6MmABX9pwFH7iKmEfvsDu3sMRW2T20ueUlC9dWBuRtDr7AH2/RLM2gph1aGppbpojwYGui
+zWYy9a9qHbaSlr4hyGbgWjJgiLNVCcnejSlRSUA226fuvE2uP02nvmFlba6qiixvkY42eTmSyn+
SLE6DZdkr1w98aU0vqILg7piOzBq5/XImwrReB+1sbfljoIujL+N7wHfOpkRYxRA5P5gNgigkYIP
vXcErCPjamwXMKubYfUWAOe7zE8eao068pBgW7sao8NmBXOVfT5UJHvbdPM3E5Dkp14h7WUbby1V
4WtQDby27BbR+oAkl6xc/rttczHJhNMEe6bihuDN+GlGD84zZpgzhd0cTIbGdtNJDcBBVTKSXBn7
Kei95ZPuXX8Q8M2Ow93F+NC9xDIaCiQ4uDyPBWCy0p2ttaQlBc+qwO49z09HyBzzM3BjWTte1W0d
jeIyvt4POWDW42tQplrPIF3yk43j0NBsn+It2G38uxTB96fHZphseaU3T3I+awEhXoMNAWKGK76e
HSMZX4n7KQDGSQVPQ6QZP+Vx8nPcNw42NoLJFI2v2Sw9l36rPVPuDKCr9OPn/ex0F7T280EsOeNy
TwzRBzhANqSAZtuNR/mYloVQAm202v0Jr+L4A7C6uJY9N4rwC1Y3R+uUfbG2AiGwon9I52TL9ykL
SLEqULomKe0+djkhxoSRdLBTM85aZk8OdKLtUCiu8FJW+NhcIdMH7bP5ilPB7KJS5Um7+nTVWlXy
vM0Psw1JY26w4UmJ2+4u/Um0tuhuUYomhlYZJFha9mB/FEmEEQ2oaV/246loID45Srfyu/NrRMhW
+vZGjPpsjknIXY5wZaFBipQjysnTNw1EFXufASU4cEgqLQjiOSCqIhOf0GGkRqe9MEOEl6cYq5IA
iwLJzPLR5UcL5BqyLir1ykGDaz84GdIihodBl1O8PzGLwcb001RFgMPYXEsy8Y9gbFUwRagaOs+7
B1d9cvpAtKvcf+BSJE7jgO36evbD3u7g2xD22b1z4JCnsqCFudU6Lx2pkuvORpb0c6nPmSSdtVdB
q3bAO0Knji7LO0bvwDMskrcm0nWGTFJ7zqv6An1GY94YI7uqB7Y45DnQuhoqrOAvxgji+wB5CPhY
b9r2QGES+/Tpz/WKHqPE3JTTRayKV6XjaJrPWvPMY5a+zJ4VnvPM5isf4K6CjnIp7DNoVkCqO89B
irH5yxIgbBL4BlTN20WSropBnkWGbRfgYgnRIHKIUwztkraCvLqFzyJ4QYuVvr0zUH09O+MVhAtB
a1/daRQGzPKEeCqf7HeMyrebGt9RLxJuExOJl+kLyvh+7mvfTeCXTCiw4Wes2TCVulI+z1XSgmf1
je8IE3tqB7AEFdyc/9KvQiz3AUnLNYWsk/ePtSmj1ypx27dSGPXeFK+RuFJbWBB9+C9YAKKOqWus
AYMw14lq8W1pFMrCfQblOhin6A5gOSWlz/to3Nw68JjxLU0Ak/ScWoPMU208iUY1cgoH9IxtXbX3
7u2B/G9WxOVasjZFfa2RIFUz0Uh9ShAYHEwGMLY+ErBRfb5M+M0Qbk45LtQ3rgjXgCut41sg/Mrr
YjNnOLcWEMqIwdoWiGhZaPPmP/j9V4W1d+UM0zdq78GexixWmf8fDySK+j2/7+TYp2R4IKR8mPfT
DpU9ppDmw7Sk+lCUo//cqmkbnGVlwQEs766n/Fnm7R9/KVz9pOBbSO4gsfZz9YpP30vOVCvVFYwL
LpM6R8SzNXmapQC38zHtB3nsaFSPSC8Ny/6kDsjLVGbSvDiVYk9vVRNU8m3YW6qhu5HX2VpmOBS5
VPbMi6f/IMyFZCeiUfZNkHjZuCS2S0Hin2r0Xg7OrPQ3QfyhpYp0PKEe7I4VzYEnNnBkw3O4GvUe
XiIzlubksrU5P+ijl1yw4LAB831lT6h85RJBsqipI4kXmsDYf9tubMBHUazHKVZIMwamAsOjTUo2
sZlok0Gq+5xeAlKJMCW+Ij2dy+GMoxdBixuljWD6M42/W/VouAAEzvZRsB9xzbE49J3pqBBdQeuL
RzK604uWzEwef1XvdCE5CXaiTt565DqxLP6Lc7xPbdwCUtGebKKGOGFH6oqQR59ghlAZfg28LJAN
NkIpL4muMAsdPPMJMj5/pIuV5VswwxnbcXqNbuteqs1aJbKS9RhCRfExYQkBNra+NwJm7z4FF3LH
5hUylI6PhzjDPG51m5tgHv87P9PlMLRbjg/krg9Bjrks8yfY5FAaH/G1WMeIB2XGnhO3HFpaqE3n
PJKz6lkIX4OvhkVqqTle6Hp0cQDKTL7/ynwIpjsz/+eWL6En0MX4OU6ZNGm3UXrSs0gxOmmyCCUz
KubiHgnuxk8T0oGJX2yHoh+CDwW5mq+4stpceZp86CQdl75Ca0TKEbNd2HHoLCz483e6YaJmkTD+
O+f63qhs79YJUpuc1qAltV6CJmwHQLT0I2KwA3NuZBUo5hbrlhH8imwBwQ+KvQAe+y+Nf6xbz77/
yW5ORausqkM94kd0MEWoE4LlDD9uXU2/sUdkYq4y3FrtgXLKbrCuBMP8iJGbfqOjS7zIHucfQH97
DcMq3ADXVv/vPm/ybNIYJOsZA7cNpEiP17DBf2cYqMqKzsWSRi4xdzCNSh7zrLfBhrvKYbkALhD1
l7g+k19pykNEjwZ4QiAihg/mFObRch2MFBUwf4OH2h+3NVk7/1/HA001394VttvWxQ/tsioC+aNY
TyyW571mwSN4osyTwrHHXGbFLtT7jUY3ff0YrYPYUzMY5aSS7+wmkFrpXAasK60c/EOdSLsJ65Ap
ne24Jmb5nyKyFHsPtxUW6fUmIz5pDPmx656jwHXV/Vf3Ohlk+mwTEnyXi+kBjEgcflMEKIKrfTWa
m6af/q5NTX05txEtBSK0Mrkr5Ilqk0GhGQE9tYtLwX0Z08wSLqL8c0pqBZimCOdD6XEo8NeolMbe
Usr+TeoWaSCpbTJvT9skcH8h3Uz0PoVrIwFy/HgtYnVVjN234N4e6TC7SjWk3+zC+nFV2dxTUNKQ
v1UemvW3LBY/qL2VDA+zDvwdgGjxqmvqKClK7GrmjVi0v4gahEfjgVmCNOnbxA1HSiO+bOBSBUtz
/2lmemVSGh7wBB/QgM5R65rOBrnY2zwV+aJSUmi0Iw90dY8szJqMMwr7/wJN3mj7jBDD39o6HyNq
Z5X7uSa1Yjp4RpUIZPADpNr8v3IcXfuzoHf1Bmlq7ntQPB6IqH2TUcL2Pv99SN6WHLs++D1f2Tth
/rxEDFNucSyA4Z9qvGXMUSI/SPtd9iIEJSW3kB0xLHsIhCaX1y6BGFtwecFDD9GzeHSfWCXSppZt
VZ+yn2VutOun4Mg1P/oel1syHWaXlLk6jlnKXhoxMuOrHQhfMnzQCa7SIvasbdwEzNURnoVNA51s
bpWOkjdB9wfTz3kEXHYJ32Q0b3ZzmbGngUr2pkqQxyjol+Q1HBLzAL4VJB/q9i44uDSTaHNXt15p
2lOiM5GiP786O7LkUbJp1FOPr/O3h8x8QzN/wp9lCUzPeKq6nx8EsbMrC09+X+mK0shkTakqeGae
okLESrihzz+LzNZ/dgZ3NbpNaU7DrbNlHgfyqJdazmzSZ+X7Y1pZgCQvzj3ALljFggnQ1qS4ONfP
l6gB82ayj7KIjBWoXHARYUYW5fOxv7hx5poDY530Fbn9hTLyoLgPrlDMmNRHDqOE5FMotm+BShpn
rh5OYQWKEskOqFLHyFJPJHv0/dCe7cYkfGkYhOurvPHR3NiY5COsgHh6/8kcht5jYV22vUStPxBf
79bpiNgXhF1r2gRljhx8ruIROyaGiRmmZbYZ4OWSRygFdPMUrfQDhV63GkXt8UGcNpjuRkWMWNzX
YAD5VlWzRWkmaKVT5zHfPqU33Jnt/b0GFDEzvKNMW/69SeI+6GwMrjasq+XEfTqUKerCKo2uTiO1
gOzrxRoGpDg0y4eclpWPH9HGetsiPVmPrpPxfnhizDXdX4VGM1NePUlixlqllQOhItxd8ekylwBM
gZgZzBc3tnQRXg4gEUnQ0/oBuBwS5jJ6dQCXcthPOBHxIrDNXM+0cH/Zy8UY+WFFjsDi81mcRDko
yEyFybsAyyimIzw5W6EM8I2mkrpB3oXy6yqchPQzWdwwCHKxbxJH0MPOigMOHO6lkNOJ+T1eGYeo
JARktTCqpAsshMX0boK6jonRyAe9dkD/t4TPMzELzrC2C7gfnQ+brVyYg5/q/ffx2OQpIHBLlt5r
CFwsLAzlgN83+jE07T+VRfJW6aNXmsSYEvzwfdB2o+sFMwXjCNPmbifJaqD6gMC01gRe+NTpLpuG
fo8ADuXebavGZ1Gvmbrl/MUT6Va1kf0sB0ybRWg01aOFUzh0AZ+SXK5qffrFpX2q/OGUmtW6SWNN
Y13xRDpDxQ6Lbv6BieM/Y5tKIR7Fu8NdRYNyL0MuXMYloDpfrJbwzD1z1xCqPH0fBK4Pxa5oZoqW
q04rhH9Cj0SfLpTIzj7VXIX8y5l3kvOm+jMOdL5otFSmsYxC+nYafU6l0XCWJ+LcTJrwv+TSHZxN
TwhkowqZbneZBYHL3dueYXgZkA3zIqhRZQ4HxRSaSoNII1yGTozUF3RiYi2UzAcf0u/xEOhAsLxN
zx0SICg5n4b5GtiQeNxDbWM+qwOPPxIt3XT1tt1pT0VJdW+4OyV0mWn3u0FYISDg97+GTNyjAt8A
xOXndZ7J7Cvyt4smsurQYWw99MYPEkXY4dKTblLaUnCBOMKZv1j9P4r+ZN3sxucs/+Y/OGLmRO2s
vsGLrTi2miS26nRHPuCaWraUhRk2Cyh3Gu1rhRWPcQgtSPoZbD3XJMOUqKZYuolgGTLr8CqslkgY
pIJrAm6Ru3yeUP11skPoeXDnJgxcXoILujF9dyhOvLvEqilCef5b2aaY7jJUn5JDr9KaEayv/Oec
1FNiCMkXh2tv2TYFnDr1w9xGTIRfHMKXQohHaKMEqEPsIoV2hlDyX5ynV+y54xxJ/BVZQl3RDZtY
OnEENmwjFtow+VmsBXp24S0rl81Ihd0xgLzb8oDMShHJQFPd0w0EPTKEpjrw/B9NJnpBICzJ8OnX
orGNNkQ+6wF0Akm+ETxM/+k6b74tRPDt2lBRWaz4OACJVstZlrOuCHvOhFIfpL8efGBVV4u4oh74
IC9eqqehMwL42bdsrtyFipYnCbOBYj1rNhwI6YforrKmJO30CXNhAfNFXxlypbQC3o+TOMnGqNJg
bUFF4q5vqRm1o/DNG+zKZhC6TA4EojNqqucNMZ8yNPrk+hR8t3oHkefMhh9w4ED6K4/vpx23M/hM
izmVkeXoJ8Dr4+a7xGmx19M6MaU5gsC8S0rGTGfPaOm1M2Nzj8RwpEF8KW/VpMr0F67a8TheDyof
m3dNg53kXa4Utbc9IXub8sXVBxd2DxGOPZXa5rUJ73VxAjaMBmj/+NA/UXtAbcA5RsM9XUUiJgEo
zzWeFTTtyLOALeue6IagFjhZZjggZaZZzjyeaU/TUYBXOvoV4qJScq/StPVyGRF8wQj2B2DpyN73
kySjUQTAeofjpFXtbzkfmcnW8TZFay5W0WmnHzcozC8FOzs6tZMH8KzCOvtIw79Lu8f0i+KzpWoX
lohyTHfdniNjUNiVNtF0QezuEeSfAeR9HYOs3Xn2iiY5vyb0BT7KSkD4bvZ9fWyg5G294mYQnz0I
g8qDglzRAtlZtRrz0IGlDk0XnWKeb0DUYSjKcDsLgRBqT1ppkJlN26LrRPHG2CuJACM3fd60fzzv
d8SX7BMBG3ABcjoWqV+Zfy/zLv53TU1/JhfpquT0A4YxOZrX9g3PJ9J8YYiLEJXWnuHSKVfc9N2b
BNiYLzdcW6ToD2p0NV+OlkLMhknJDEfFvUs2HeDhJaSZQNP3gPKBqbFVhXoAjcGa3zb1AKgFobQp
6QGIPM7ujLTmK3/aS55EGm/mVtE4+SX1FzX3j9Fb+Q0HkxLT5ZU0wBm2vYm2FZJ4snPdv6Ybesqb
sAY+xbrS0VEhOmJyTuN+vGU1WwNzdvDSihaCMGP8ozIlykrtMZHeyrQ0q8VXXI4LdK+j2tdkESPR
UQmQQUjGR4gib6I/Mozt2RAW66Gy3RbJDhRzU+evCGX59lVQFun2YdD6hn07rlM8PGxztpzy2gdc
KDdi9sCMntDat9rB7wqFufF5C46/MzWL8zm9rZQGfP/4el6aQBzjU/dTDK/4U64inHDnhrI9Bxy4
vs3tMjbCtEGHv3Io/dRtvTI45/B2D766vAsUmFdEEIIhiDanAfcquMW53O1NfytIRXpAXwYYKmUz
7KmlUbxjUYpNBd/OF6Bk15MDTzOdPv6sIp01b59BXJScwnoUrOoAsemAMvUWa61tsssDA78f32hF
cKLSXivdbS6Vl6K9S8+eIWWcweZ1FRTQK1YznOrSnso8JoVddMk7mCIXp/anQTQSfxZ4e4Ys7G4A
UK4BYDFF5UV/k5vaUaQDddZrt5mEuYRT9sQtF+K5V6lAU+Ma5vtafqmo6Cxmfvhve0X6KQ+3JEq7
oTu9ewRjbx9sxTt4MF5ZR609+Bv6L2IGRm2bkyprJVVHV7WMraTYY31LrdJ/tD9Pu5T5S+yUrp7t
1qP8QN2D8AU+ThH2wMZGrZpMZEi90p2lIzdNKTBmej55zA9gMe6URgbApl7zOL9OIJ+exSxu7elW
ssiKZ2t+eCrsL8WGbbdYHfzRn0BfLX9PXDFxMvLM7240gImtC/1elpx/P0DvZAMJV0X5pmXCj4oF
q4SSh2IMmymZVHNyHM6HMaJSbINcOXMLeFJwVt5heJS/MKnYfy0/c/ea6dyVcuDDG+FA6FHjhtRp
JPn/eqUmbuaCRJQMiKhgG9JVp5xnqMnojc0ocg9znkckMVVSNpxMgrSETiaglqSsOSg3JIvlVMfu
Kf20Ydu8ysxf2PmdN6fnoGkj3FdPc9ZR0ekge5ci9diQxvMcClEun2r6Jy4OlqkCK4Wox2qr99iu
sTHeylYzIzE0yQ5P+MU/6gR6MyFJYCD4SigafVI6MdGCzf2Dg3M/xFRCZvcpEyw3gihm9plb6zq/
Y8BSemjSuYE4I0wtSx5n+mvZLGms4NbyLanA/LV0o59rqENswGX2x76wYXxc9lnU9TfokeEkdj90
0NXbH4gVlt+HkeCqrcgczKIAlqwLvoD1FwUMooAi0OCe/HKE207V74nOmR2wVRSxp/Awc5Ff01GT
kK94mqv2plO1Rv9NStnYRFXk7e/8aqfP4lEgiHpIl9qAhPgmNZ+T9pC1P9yGkBi1TbKeOc8AqVR3
q3PlztNIqAnQzos088xVdy+SobqDtFMI9N1mYkioB+InleCvWXlXvi8oJUiLi7Cl36uHoRn9p3Xs
wXKtLdvqHy04R6B/cN6lxgMADmKss+27u8J16D6d637UPjCSIdDXizb9v4cJ6do/qLIXgi5DPzwR
PJ7E9aiRJFskHyc6HrK5Laqi81nVit6R5h9or+XPzLq0mh7NzUPfoc+JDxdCFoLDg6AnDlr+Z3RG
aHOxizL2o33Qea61hl7Ah9H/V3ZicIKFd5KLVB140n2+qnQmLLrJv/dr4BjMUoNKJpzbBXKscK8E
g3rgvgRaUCwH929VLz3KnfYJBfqupWoej5PGIqSMcGLiTO3B9Coii5VTi+9t30xB7harKb8xw0xM
rnnqxQ0h68Msvax5WnCWhDn5hnDhLB4IDDOh0eBcC7uwJuDuN1yChS2yZA1CdLqRvTANmQYNus30
WYy7AIqas2cFeRd4ivC7l9LlYRgKazYRuNK6QyHHmZuPScDkqinXUW4PP8rDGTQiD1YXt0QeSOEh
38C1lfRuh7N/KOz+94/2Od7mPW4xKMYVDtYsUkXy6gdxkr3JxLmUGMwEMbNKuglGrjwPRiBNS2sC
I/qs7VEZUFNAoHydmLlyYdj7w5lnhlo/fgDDex7RBa6BTyGagq//4PZgKzrE9SoZUloEPu7sFZAY
2TYYp4nrl4z4I//rwF2q0ca930pM5q1zkksaUN0hZlfBnSGs1GzvpY3zWSZq+EY2J4oFhsTW6V6W
R/76di2moMyT1UaTIXdNp1QYlFo0oKGXNWkG8IInZFQiL9yT//j9n3Ojs2IWIcZyypdgd93GiU8R
gJs8fhu9HPn9FJ4EV20cgcrxgePoaAZXvZwcQmumLGp3jwCkVuzg/4eJs+ITcWK5LHyUYofOL1Xz
oK3HF4eyuDfnI5EaQ+6Z+c8as967JByhAcj7T2fQsgJ1DXlE02wO/oOYISl4f+ticdCUbCUcqX0k
gpNuWRKy7RPpTftMX4FX5RhDG/xPwTQt+K8XU9blaxD0nA6770Sar7j3t/OGQQMzxpu3yuedraSQ
WBvka6ClkxeYcrgpyLXG5GHg0Wj+r9FljGiP02AMRRHVfCTmpZ4/a4UAH01Px4RKDjo5i/w/KNip
xG3pom0AveAEYWTFNj+uz5WmGAH6t/LuZT9Cl6xFZX98YtCrn5kfms7O6j8o2BmozCrXUJz0MKRG
7/OHmYJT3HAMzUNb7ONXC/rFoDazSSWzqZA61UlDdJZzu1Y2j0mCid2Eg4eXIm9r32+zYCxCAGRx
KnMfpX0rx38CWQMdknZsBN49LDfj5Oz5HQ3dy4ivroPs3iTK5WhCzuSV8FUHY7HINZacVTOGJ/Dy
cRGqEGiwYHvIch+hQg8+cu8pN3ZVf9WXMi9PfDAR38m853QhqVLH1Ph7wYpJJQ8r9KBjh86RNEDQ
QJTaIcnMvbDXQhBneFYP8QEzh+4kEqqrBBWnlt5ncQkFQIGOXSXT2Fj6t8315zUArWcRyD2fEiS1
eC8zLZwoO3SFXdCyQHjx8KER6vsl3cdJALbk3fZVGC6SqDe5NzaaDTpScXBtPQ5+LUczg/RSaTyH
BiUTXMAMNV2LRwqNA3StGCUKlRWfgUJUyH81qqg0hDFCqbT63yu9QpAqABmNTUDHikZoHbiCx2pf
iuy/F+xEaK6mRdJLnEOGFfPb4Ft+QiifC3zQhXXPCI2q5M90ICAanyc0xiD3i8k/932gu7e04DM2
5N7IXiv79++uz2oNtLC+aAslJpiYcqscgFuzt8n/dDPEscb1qUB1FjegkdJcmqw6RyjJIMdGk0Sc
/o9RUN7N2AcLzw8qlWdtvNch57S+bN+exqU76qPeaEDeG0Yg0DeTgCrRmHhaYt+P3oZijBeQBI/J
qf7C2cIM719ff/8SBYrtKJN57z2ug1896HlBG/EAZfgS3H1z93AE2EV1movseni/rdzETsS7VlYs
dawOvXwoFHOEe3hJxssp0pGijveV6cZxxhpsXhLUlhKZfXr5koDIUGHetkcVjk4FMak7YoN1aPb5
r3Gdu7XShmL/5yKW90yfo4ewOGFktFV0hwpWrcMUJJ3ZHLr8jdBb5G56Ma0VYRyqCXkieIgB69/b
4GL1/e5DPDbFZQktwpicExBVIIQJCib4Ab+8Dz1TfAyrY6Iw16XBUgk3MbSsijiMnvGIkrrzbsQn
bylqAZ7NS/ZbfeRzOKcPrr5kht+qmQdQGvPAEFqrFf2mjr2LL5vJti157FpQhC2PSp0+fM8cHBeB
Kra8kgLOa3n1/3Va0pRw5Wke7KKb31uUR62lM0KXTb0gaqRmwZeNIDcUyeAWT/Qm+AcjY8VumYsZ
R+qXW9/Xn89jKMTOv5hOOiDw+/82sgCWCeZNitn9n6bd6GGFLL4lZKtpHkFv1PJAOQECxZLODvGG
jQ/Pz9WoCdsRSw4hOfp2UsfF6h179ET8in/8IkaslWpWGirC6COda0EdtiFQTo/OiB97eV0r7fv+
H5Hp22NKKLnbY86Jts4tfJ/j1o5QQfuf5HQu/m8i5aB0OQcJCYaZcC2/r7Z2saCdZ57l/3OzWbFX
ELtheoQ9h0s8a2vnCMyDQniThWZYM93XLqxCmXz3wRxbcXvJkbqi6ayDNxHj6Ck309S6s4TXBzDo
2h/Z9m3qSAJmPGQwugT0camCJ+jR5w4AyaBKjS8rrPjq4fJ3S0lqYK7rfjEc2dCtDi97WNsKGuxa
HDxCWI5P1mCVUmUFunfwSvZxqXxUWJVSMCUDOsgkRxM0zMPcXmJcW8G6i1JlVujSqcGSTD8PcJHV
c6EwbnS+IFONuRY0oMm+BVJP3C2qJTjLtcfRrI2gZkTlig8Roj+IZfYuuDNCze0YVpTJ9YvercTw
xCw+Zfita2MAujIo6ss+YpxWU5y4MojLQxjJsqzvvKRgf0QPG8CMPyouPYrIx17rtEHw3z2y0dOP
SxU1iFvPp+Vz2AIIygrNOn0J1WiMrHf0IC6JlN15uC+p3sIdwa9otlfzQnIlGXhHEd0P9im3qVzS
vvx9QKU24AhQ/ageyuf0elB5ztP1uDy2Eb4tb1EMVk6M1Y0V+epfVvxwXwmdCl9UALzT5Fh4YmTW
6dtAsxaaJsnXd1H7w6wMxx3ehqTrR8qQ1am+e+wd99tvxJ4Xjo8gOxtk0mXWlAGdbTwuo0stKAzg
YO7IadtYgo97cJqMR5jpOSgN59W6AWSeic4+7DNECiQ/Pd7iiInGSXT6k14N+pRcfFnYj35fnlBM
FMhprlgeFisFKNIWwTMu0RvyeWVItjkW/0UL+oAoAo4UG7qHv2fsMO1LVYEnEoVnOD8ty2pwwal4
JJvnIo2F4/j7cl+4qu84O/ikDhRANO6ykhfV00aKN+cxNFKUIp1+TIDvewrV9OAtSX3Mdu+BiQLl
kbJMQ1jISJNOvlYwh/q85PsJ9vO7D2WkUW8x7xmgf95/FDjP91ljfg/aJMWvrQtuV8pI23l89eGT
UN9Bfr/HX8wfCcUgV8Pzq07fWw+TvioXBcs0N1SvVg8NNqj6QEY5jHIuZPvtlumCHABKgwF0CSeB
cK70ZJ7r0muKebIqgOKzL3n01TXQlEJNdDSFOUoqUuJimqSixxIdvwhsyhMaymWF3vLQVKafRP8O
klub7xCMUb2WWZtekzGKZJOx4iWcSo4d737lUK0xpMSy/obbFcduyYR4+bjjNhbLbmnFpdE6gu9N
Q2S9C3/sWy/Nwa+Qd6qemZgEiMKxYP8dzJYjwSgmLobs4D1vLCS71mYhz3/tJEZYAxpMbq3NFMWA
n2HkA6SQJg7FWgfUt9KNKupHnfjzjo/c0JkAbbfdFXHX8knzmrrW+cQmTph4+QPngb8xEdiIpypP
WGW8USC47D0AIh4X7zxC6Mxrqp1aTw1jH7iPgFBYlnqelozpHpoHkshp+pQujip9WeVuuO1qX9Ap
sR050nbYj6TX0p5qf3ip0HBTnvvlvjO0arnWNTSaRyeDw/CTd9FZ+ie2C/jNrx4hmvPb0f7fngjl
ni4XmBa7Mt9U9nDvRkAbWX89s+CfwM5CWhVAAfrS8nRD7tr15bJUUVQIUg9q+2FRNo7Uc0XiOFsq
afu7llzbXQ/2NXLBBwIxT6sFyoGQfGobHQtoC/2Sz7Rta8E+GGf0s5PSKoZ1lr+UJ2yXHydIoEKp
vDwk/FMfI+2Jbx7koV8bUniJhRqX1s8H6uigGTr5U4YVLcWED7tIQptZ3+33WFrL/u0r5aec7x3m
Nm1vmz3ToZ+Goor5VZdWL1NwjaDqW9yeyhzEo7mkW0B7AaAI3KW+dpZT5wYwN48uv3MwUiPWCn94
0IPyx443iYSseiaHSzakDY6Nw2z8yd+wRJsKAdpofHBlJ9bxoWUvVKA3fr7ypNTnEGcPOSOdIQeR
kdilssXvqRUtMoEawglGVCx91yb4Bfj79u52du/zHB4yWlN2ecogpQvt9TSIQCzamtzJx5Jj6hSN
Vc4s3oERCjxgl7NzAhOFTfihc4bJDsLWwyNRtShPodG0OPgNRn2CUm9vtKxqOkPOCypEdqvr1pIF
QdvY0b3L8uJIbkfDxinppBeEVzNc8das/pCT8fEXpeEXz3aLdNANppS+S2tf15c3EeFhMqDFafrQ
KrgnXjplMxV45B7wefOOEX7h1FJYue4K5hdQHKJG42PW2ei47MPH5RQVrzn+U69w6l88x9oXRYl/
nzs0J3t+FFj5kHl+xAdYuKBCuhOqpG85FfKZRfhHNF+8feNQ8K2raQUaWFGmX0vDBQ3CvuMNV8Ti
fymS45lNwYKSfq7BGAt+oC8mCPN2T6EaqzpW/2qtpxsNrJUV+7DYQGoskoN9Y+HXX2uV0X90xJJ1
wz7RtQqipUdJ8Ti6ZqQDfYfBME8RyRdijA9VcUAp0Ie4UcWNDtwLK1xJoU/Sto5rLnruXzuMCjKC
p5ngN7Eu3Rfd6z7NX3O1QAstep2PvezXNqxy2Ek5Q4evKsl5k6Esh3C0NDDgPvI/MxPb3wM+/NnD
jLdN1VJOSGdASuNtYuyr+/SAGYSX+dBKCn7uw6hTUnvUf5MRbzCfzrOtK0Be1RDOAKJ7RK7pLBkk
vN2iWC1yy9MhNuy1PpR3OIkLVuFxXvov2mniLQ51Jcjl7ir5t6D7u9LRu/5HGs779mAwQXRaPnd2
C5ub+45GtndfYmMP9S7sd3PE+7+MP87qavIM+KGsFPQ9QtHd/cWk0Z1IHU4sM3Q2np9VLIgyOwCZ
zYHX7g14CMTChcvOhvE1GKi6qwmWMY8+8wli1x9nMCjNUvQbAxRJieGrPK03A9NeM7zYAbxfj7D4
aJj+7a5AH+My2LWhfHca2CtcDJcF7ikdDMrNedW3Ohd8pO5H99ZtYdL2W6vZnVMr3goTYL3kzK22
Cw923aocFbJ3LBB53FxUHHn4ORV+Z6fkTvKGEaQKGh2JA9usB1ICGFUK4zTBHHTh5YOQUFfChLyw
NnHu2BTwowlEMuuJ71cEJ2u4hodphKZnsc3o3D2x0ayii4r3J5wvtGHGCCMxCygIpnuJcqDyneBT
KytllkmrB62GkaoNESILh0ITvghgyiBdhrXlyWzyWsx59A9N/fAItahiT+2o80ZcvZcxBMx5oqOv
dMVmntCQzNO+uRlqQZw6SlzZhT9jLpZjrpinPQUgTTB4FK9unAsdLAoq7D8jLFVT+01gXtz1vrAG
zxZww4X6Cgfkxy1HJsuKmceiXFH3A+SjYkBNeADKGH7jUipDd3p/aMpi+pOAtjPIN4NAsvN0bH9Z
AuMGbIID9Il/XGdJfdScL7hf1FKCtieGw5KMEd90a3oAB39q0VtTXH6ci3vgRbP4gfhVHDgwfglm
Gc3eCzodoLjlDbc68PTA4e+XxTQoqwrtYAuC9H+ot1ERAQHK2tV/nEDz/gsg3vAzjBC2PrWtkmfW
ytX3WyGHWVk8v1YUdKTGaqq+SHM3aHj4jRiHKkxeYnD4bY/TVH04y0QS6i+xedktCBnxFL3h+PWn
0HDZQfiovQAkLQSZY+njvM2ar4e3WS27YmcdtYJ+Nh+i3eOegMfVoxSwmd+GQ6G4EeCWxVk4CkhT
kLJjG/oqdSz6SXxB12TIlIba5tocmje0+4jOZkE0pm3d34Bgs0NgFYKQJizkMUnrdBeueWg20/2Y
vUpIg6R9v9oCNoq36Kc+EhBMKT37T49Dss9awCLeGvtq6ytoZDbFqXOHDpzbK3pZ3PnLzuImOm+O
qrW2lmTdMmgdyLof49MVxiZKURjTuVGYSBzQpsgdHVR5Aa92k3x3Ana5vIPQO0alqrZ2QffhE7mu
W8vVJMw4FYSkdXktKtpR00EuykdvZXws1qJCkBpxP68y0VOM0P0osX1cW4z+MfjakS0AzpZFqH1M
JjXvopqDODqNsHopk/T+tkOWYBV6O20mEQBfeHQUvaBDycxKjF5lUs80ahuadwzqxGB3j9YdiXzn
9RHnwAXyrqZeXKzPorl0jNi1K25f0UA738sPy7NFzMXk5gEOwOAfUg/bQdHEHsatw/eruZe8ivIY
B+TqjH/8N3AT40Ki9p1Pp/45zUS2NgH8WcxH98KKjkxwy8mZu8r6ey7Fa7YCMO4kR3mOxY/LUtnK
pTSryVs6/oyjGjDI8NW7S17fG8IAewZs322uKtF5sv8LBP8w+jArGWzFiSek8CtFwoZCYtKCpAwr
g8op57XETGPtDE/X57cgdP2D+RoMXoOLA2NGHgscIiD79yskhSlt9M84H0X2t4icnVuzRxZzvSxT
fRR7A5GFMEYuPcOVoBP7kLotn0aAOHa5KAEIdgtyMrcZT4nEBfMDbTgsFBCc3KieTgJiefU9vU3l
4Fai/gPz8VVnGanIdbKrDvzA4faZoCn/NCRGkKJghw3P+QEjGMR9FKWTLMsUJMkvxK4Lk1xAW5j9
HB/eBzDNcDtqD0k1fggJfnWozNZNFOMWFDumZGCe3lxo3w5qZtxRgpZOzIV775WC1DbzVbsw3MCx
jrKOq1BqEUD0g0ikVhkj058aMtNKDdjEl22RR+NfFMakccsRLrGFwYCE6vgKDpuWO9xDx35n862P
ZpRQUnkcsVv1E26OsMNefloJ1KOt0Mh6OoEZ+CpFjCy4QRqgk0eM5l0igMSZJOA9j1cLMQLuuTPu
2JVFppyjWLCV1gNQYzgqRkd82aUW9O1uL+G3v9RL6ceNBPpHzR/gqj6yhOV8MaARIDPYTtfC69tB
TvVoIGAoScJ3tkVIQ7x7V0dpL8Aq20XJQZtz5kszbGYMum76+79dKgEMICfA0YgazQU6oAt/lBBE
l26Ii3QQe4otvr3JgkVrY1S5/xl6dfTE68QMqPsA3+Sh6o5o9igIREcPyFbyn+O17FcFTcbuXCX0
3E5T50Bh7OjcHo1fIsc/NKNKwG+0oBeKnpRGFVFcZreTXXb+0si6HxMIDIIV+jvJYpbtc8gTkq2U
t5gNHYiv9v9lHhwM+QyLoYkY9v4Q/vd5iehlwAt826imHLO2kmdzR13yHddCiZTLDYjzKWUjrdKW
ySEB+v85ByyuFlyFrFdh+xi1nM+77pMeir2iCjAmCeHLiPtzC57nhiAXlwbdUbAa4n+3dZ+kUi6n
okLT6q90lz+Zjm+90y8hYGiIIcp7Vy9nRBDlWqyyEJTIXj7UennQJ4HVyyONtaPkD93foSYYsAR9
l16eQo07lai38oDDIp/SNDsdYBAWnuywWMbb6jnW6ay8R10/V8JiXVvuhLWxCjrbL76FFtdrPMPW
SBcq2IteE4yyYusytUVCRN6Pt5DoLLvXfnOASlW8YW8ptaOxjcy+Pb0umug0wGSQOm/5MNjAFHPZ
UQrUuyf9LybewrR9fLyuHILr8ViOfRvwncqZWeMlXGtpul3IaWe5MMQ+ojmJA0uAqSgvyDKiF34D
0azMa2DZbZFhUmlOlnFrQraWtDjxJwOGYV19N/Btvb8NxdlGA9OpFRJxrUwvb0kWpHtP1RPeW/Zk
Xw7yao2KJzQwU+HsirmS5FGN29fP/+QQodscpXL34eBp9JPuk1GCqkCfsdeOGNTIUfjMrC+8anzm
JkdvS9uStQ+bgwo+EbT1IQVoji/WS28XiDK+p2hT3cN6nPP9dz4elr6Tazpb7XfogsqK+xvY1ImM
emGA+0BQqaQhSshewCYMYEZCM8hrdo0X2Yw7a5yVMPZ2vR3qeQM+08EZBozPeW0IBGkk3/Tot+4h
wiDV54+yzfMPQYfdCcJCJt3tX6zteklx5KSLStv/9Vg2rL8mGNjCTcEbpwl0kzAGyJCTRKJqOs0j
EpikmLjZwdUy3Lj7Lh4m/Y2yQTI0AKUhmuAp0SMZopfXX4zVFNuzG05+OxTKoPGiLpkmlaSh0YXH
m8jJJLwbFdClFgUgOZ7aRD+qZZC+McTP2TG/Pedw0m22LEQbIte9fAv5OBTCiHPMPHmcUSVXtd2P
z6V7+qokzBMhlm0LRcSnYgW9JvDghImlb1IWQRhwxo6BfPiJ5hbMjmg3w5gSKocHkuDfaDHcUxjv
ROLaKOsn37THrJtIdY+faZXqg4uu57k752l585XINR/OfLV2cyXK2E6DXUT0vlMLPalzxN1ZlsOM
JfWCU5s5ygIONGURnJszBGeczCwc/OcH1qZmXymDODlWzy+qNcaIfFX/EGTrwdeYDSYuTz91DX0Q
g8n3EX9EIkbZ0ap4+THHXZrDS3+O7qecLW6LkJrbi9SOiBd24TqcVaDyjrOwdKuHO1RnXeU6USsP
NOKN2AHavG4PGWZbSZurA3D0nKerguyHylIyE0rbhJyEfk7c4TXvktBeaLHd7sYOk0EHfw9d8lPx
LNuyTpiIpky1VMrhexNVwyxbZDBLJZQETPxHN+F1AF6Y45xUfEPbKN4xYByrnKRaNN/Fk62dk7W6
tMkXLoqDvBr4D/HcrBNVmc2dHgR2trnLKHblWKCPEDQ6oPAbrRfxVESosD3EdvmNIzSq2luFORpX
GEMzy/XrMUyhTocGKIckJ2dOunGaNKuBiqDZgb3NVeIHt21ji3Uaaeru2Id+5YmG+4PmAv/MH1gE
+7g8EM7+SNBW2P2TJftdSlw9Xp1d8Jza/9ad6eC32RAd/j6qNcruAPUoAMHy1eDl096O5Bl+AYBq
ogevFJWkRMQ55hqxeNttVwzOq3a9smyjBxZbTyNnTkd/oDfdbpqlQErpVc7RDO6sQj2JTF9U1gGh
52hXncIVASGP1NUR/ol/IZI6uNHy8AWosbeHHmEL2XqQut0V5EjANoQOUSYNiJI5yuB50sBsVeEE
UmDK4v36k9x5UQm+Tp60VMj/CLpS8dzTu/lsmfpAPV5BX13kz+HMrm17x+B8pfiv7XZKSi6KRg3M
LsyIezndwY2lhhAXWRNcKbZYhppaMG8OiwPAtfF/TMHYXim1LxNd64jT6ZPfabYyHSAljfQU6KdJ
Zlf0TEsKpGigeaWrMgb6hnfhCUSnYVWatm3dXGkS/E31JWHFIRSW9JWCdhnIL6Iw8vP13ecuBFOZ
Bo9WxWnEkIKU6TiKeDuJajCC3IlZ09Sh59BlV2v9E2o+hoqEtvSg+RfFAvbkStRooLtjRf7r1dx4
Fm5A/dNPkXYVwgvVu+Qaqlag5dcEBsOqI8YYHshK1kGnDxIJZ8iGCRgTzwpZ1C/z7r9nG6hAz3Jz
5k7amQ0yunjvFSD3Z9ghmoaIuGmJa4AinjuoxcsQLJgQGbUKhm+BJmqD7HsnIHAZCixem/1YvxDc
CXed8AeWHoFk1pBpav7sNy4tnW9VDmSfei26mJsHSEh6afT1EfKpjjDIUrKU2yT3BLGHgEDrC4vT
8NjT5ZAo3qj4S8NAOzC2aWp/n8RmO6Lis/C1Og4hCeCSp4BnBtRNXGEcon0nscKwMyF4NLKJzShN
zsAQ0bgmm5WJTeXhpdXwByoKV1KckJDBAho4NEF+hFUrpiOUVcxwhqOjCGv/NsS5BSLOFgXKW4ZY
B3OEL7QTg0GCt/SfaE2leu0yKHZInTEDdZmqx0bPyKDzJcQRQUp8M45KekRN1aiP37VldHco/2DY
XG6GdvE/mPSxzfwQIb1yLIZFm2YU0ULIB1h10VcXsMyAPxGvd9mGB4e4b0z9RvDnocNYN8b7QAa/
i4Tg82yWIyWUeJbZdkxS0pIajuqw1KrQ0N2Fb41jFT17iev/rYPk/yv4mJaWjtFYa/axXykmRsWa
RQUc3SgJE6PphQoaasqIC/uWBAtPGj1LwowJZ197Grrpr6R7ol4ZAoc9hNkgidX421f+igC3bbwS
oXY43ldZfiu+BNeUK2eeTvcxgEHMVj5tpx8hDaUr14/2woWhaH+JeqmnE8SOMJNxG3Lqax9c+hCW
iIUSM+0iSlkPf7g8CD1GAaZl52Utmb7mmWB6letFYugB0iXZxLbTHsdEC7CCUnf7o6yGUUmJ3HZx
xY3DaZMkatS+00bC8Z5X4sKuIPTjXK3GBm7t1/ot/3FaT0l95QhxlgKGJ9hMVb5XcJtD22SuP5K5
SaXCKpIsNBE2G3Ec/f9+1tXbbCDAp9cHNVav/UGxpT9gCa5VFpXXjDDLYXRm/kw2CtJdv1AZ6kjm
lSQH3Q45hrsnEycsSXXNV0NtKAmHsfiH947EUMXPU3W66wS/wUWeLT+g1MLTDC5e0tpFalPtb8JU
s+fzLd8ZiltalgrGbiuDTJxbExnTmpXz1qoCPa7gxNHqiUMfqtnuo5m9dS/1qe9ZJx+OLbUaS6IT
6ubHrGQ3PpMJfNE7KlwAnLbxK4f8rDinLx8B83cMf2fyzKKY15w2Hh34IAsF6Al82cTrespNlgQv
jlSWSJJJO21h50rvv45LlAWdIoEyZl6qBBTpfYDMjm5uXOktixXkrZw9SxW5Ch/oZkbIRnEkOMUZ
QfCG3UZ7nr38WC0P1x08lqna9V7y0cl6Bseo91ywqddi/EBKDUj7Ui1VGFPYEUoPwcwHTbYojtCx
Cip6PYIbUAHSTbTM0pcAw2z4IeOqLgQiCyK2im/GOlW14hKwD0aYJziG/XeNdrIh9gLWy/0Hu3Om
i7Zm4/dePoFUPiexr39SVkrl6wdLzVl/dFuS4AnPGW8kgLzB6qElJPM+6wP7QhEKAw/h2M1yFX5/
rHQ2bL8jK/4RGcnELxYe8my1GYBJUovMgiq1a2QDVhwbZfR/CNd65a5++hMARHLBQdJyLYCLM2NJ
iu1yAyajhq3EIRE489SM4yUU6MqfbE7OJM3iYScTzs9Xa8rkWubGAPGS6Fra5mBJNDP6F4lu/Rqk
jN8KcreWnZDZ8bJNj5ka9kSnVc8mpbnlxjOPAx9NJK6/jv/U/7gxJnhxtkN0aBcSHUIPV4MhHvDY
+DyewwGg+XLpLI9TgGTCLHOmd6pLitKbjg3K9/WvWKy/MadwdHK4PuCkFq9J5qO/GN4a40sRO+NB
AqNaru4ZqlpEx/zfk6ObAYKg8IA6vFQcftxLtFwp9FSsvVwIhMNgTmigKgD/skDjyHusCKwRt7km
JUv9dlPt5jsjc9rP4XS9fQ0VbWovUEWX6JbS8UCh6WJbIxEhDx4p5u0HbT286EbUTvThSpoVrxmW
fKWFD67O07DWSkzBMQ/ZU3WQL7O4siXCTuhhx3/fPfGxG1H05v9oNdgypFLNDoIY2ZxCjKKeMm2b
wa/GKojjE8mjBcwQnpokWnNiF40QWlq6LR3BvcTX4ULxOU5AUaNneU4vUDcQQz6/0TDKk6a3NGoF
gTqtiYDOs9X8FSP3wNUJV41YTraQwadhya2OqDIMSlA+ENEuV91UJpNO9ACyRD2+Ih6rurnywK0n
HqsdeEW+xQEvc0aMgrN4zskBJEo8depo8++Wp4OrMeJR5bO53eNtX9sZt9bdmPXS8Fmw+YEnazLR
w6hyPUvp5Y28tidADmTdIn1mFH6vnmM6sNkhtVqHT15XKv15+YcJLWO+BUsLcRujBvmlaTv3H8jR
WZUnXdhsLqCWN0ygwsLvj9eIOGAmNB4V8mnZewSc5aVTVKASHCC2fp1jifDjFa8sqH9cl36Wa7yM
9UrpUkh5tQTyH1v6TTEo7CplO7ylsPkKXnpEWYZEc1e5airqUGf6rElBAOuK7+8w4vHBKG5C9hDx
0kGBCKPy6cf426GXCUsdjxYMWXsmGacf7kM7AWDkvLMMewJwRX3cwCay6p6HmYt5vmPXu9W06Ph8
0WATwYHG6+0Gd9wlk1Qg4ElJQJgKefLeqnouVd4NkR1wVmIyMVaT/i9Dmchvj8CfhcKqrTAbZ44Y
XmZcOxEemhVeC6j7eSfRuU3oxVPaXgcSV2lmzVFpHUZwNMii+edODPxKAnOaQAZaVMyqnNLD15lf
5ItAr7hj4HjEYhCr37Wdltjij3l4dPzo1ib9eTx94tTHjTKZ2Yc/f5pI0ey1gnriiGquBNDeQvkP
dIMrApMKXZrRC40x5+xGip/8fzAQkCmTG04BdTjLX4JTm2PQ+MFmBO15SiZMZ4CF2qzBE2VkajP2
pyI9CWIcQKyODHQc+NfL3C/iyyGRvu87t3JPYheqdIDkzUHAhS/A3/Ap5MU6Xrz2xRz9/ajO0/Rp
qk3lAxydInZ5A2JFSMsfsLE/YrHvAJP9895htdVKQVNQQPiSd1h0eVgGqSEo3TTZhtwrbuavlYyp
fSobjXG+zz6Tr9UMUerKNjl/TUC8Su+LCdH8tEEwPcMadyvSuX5QmYiYbHvpwX9MGB1V113Hb0z7
NxKElgdDU0nrrawxdL4G/rK4AfQjm1F2AEY1fx+hWZLXjwtjsuvN2eRj60Vnmc6w4dspzmOJdFPM
ODypcII9/kYgazQAtn/P3MCkLHOL8NDk9382zIMN2YX8Nr3Z1DpMX3FwjricfUSSbMjW6cGrYCGI
Mlh9H80JvsqdK+TgJzsvDkGGNzLPVbuAWwIZPnqy3V0PHoY+dJJLzsVP3D0LNsIYuQ1jPxsPDpZ6
L1r3wjYOM2evk8iSDdp72HROOHjFr77tAlOwf6PE4eEEMt0E7F+5+npHvFLRPwZBlKEq1r2k0dgQ
a84IJ0ft38YKXPlb+8csPhcEZ3sR0fxQqsMtB88by7/MOnvNbA+cCyucWwSuH/U34eF+j76FRT8d
TC1I9LdruBgBPtv9lfJP8y6V5EcF7bIvVrNwnw7TWMx6buBca+x4oKl3hWxr3SznbreSqnoeBE9j
txRRDS0Gkp9DDbKPR8MUERZBJmPwciqeMXrIXqJMeAPWb1nIjqRY7WdcF9cYeax0JLrEod7olaAh
jQmo5mDgSbgiYQivnyaaSpu6SVtL5T8n/aU6HNqqLWZPHKPMbHAhSNY45/lpw517I4rO79rYkxlf
o8i/3Ou8e2RhAv0Um5zx0shjoih470UOZ/Joydn+1LFXwiihgsAKQVjhe/iH9OlBtA942hCYiUHF
oLDRJpt4m6v3e0qAKQb/3TExw8ud73HBvnRB5CjeB6MfasNNG+yaslobPomHNhBnx1vpQLxFJGWw
xcGenm5xnsNOz6I95ScQz7JcSngdxDEx1DKE5S7ubh1fkc8dLWvkZvzu1sjs92xj/Cd4WNs7uHbN
Yl2B1vqNQCB0PGT+Ta7PSpmJ/URxPhJsa+xctr9ERmbhpBNWi33z0aekU0Repl4OJkCM+1v0GAwp
TDwCEpAFceI5zIdmGhBwnWLzUrOaG8SKTnZUZd1bZEu8svuDKZWwURyOckFKd9US/trh4Nc/IJ7q
3FGGZis3AVgabi5wDBNC/GXZ4TjDIl3rZRhgyqwP5+JF5rM/VJTIXkJnzV4b8Sut7xYEEDZbkWjt
ywV+HAQmVvl7cLc1kw10ioyP4v0h130Oy+5RTmycHb/555It63SL1IWYGD9tzQ01cb5w9rqDoXsH
PcejJSvlrSqRsSS9Kz2wdT7ywzCHwTJ3hcMqxHExA/aRVCa9Y1lBjGUhqIaRHG6neBWHXlA+fDjj
Chm18o6j1thU4ttm2EuTMP4LmQGV0SV9hJY3MtWD3YkMGEZI0Ug8k+19ojNETOJlgUuztj1dyxiw
J50N6DZXwqi1AL2uIwyrzysJko1hpMhqK2MxCqYpx47ZIXEj/JLkWgphFtQh99ke9zu079k8Bxtg
41TEZN4CXhnhKXK5oWql5zNcZx1Tdknxye8o2nY9OqS3I2qf1yTkel28SdooW85AWFZwQNBS3P1x
RYU25UEo0Vnu0xnVjWu6soi/CUeJDIkMyCk8PlwSYJJaAqDPPZYgrKKqe70spIseNGD1X7Ge3lR9
pScRcKXdujHmS1TpSAm/3PUZleqEBmFgcNBbw8OdL6eqQUfoKoiPwrDFUWWyppxeGOG7qnIhsqiB
MTgF+Vp43WQjeePXxjBtPExE9WiUmqytsczqC3ptGOumnMevy5TLCdw5w1/Z7q41E0yAfyN0U6qq
SvofQ3s92HOpqIk22/i8Sks+TdxvJovQQ+qttq4OldOI9fkH0Ev3E+9cXTJs4TCPVoKY75TMKlw/
bCkYmXt8qThfD1RbbdARQpkbS3S26j3KU00tSICKPxa7EqmivRqBEEDFM3srfdtBOUMi1KDF4GVB
fWyk3QdqjWzh2oYbNUMbwWS6r43pCAVMhhPXJVA9PjFRanK98fYi9hEP2TRBNt2thkAv2ML19kvO
AzvkbxZbelk1umL3ivNIGsWftl9b+jlgZMa7cWyyS4QUFPvd4Uiis8q8EE/7zKcMn+CJZtdbGneY
q55YMtp43dU7i7ZIHHCPeWHsLyS3MCOBK5HCM3g17534VXfG0RNWJvhFvmFWiBOD+ihgb/lca883
BZo5ncY6nMCjkmcWtDdh1PONsZ/Nyac3mUEGkkaPkYpQ34bl5LxG4HEE20DMDch4oSrMmlg4bpvd
4c0mNpA1paF1L2ArYRtl3tCFLQ6srzTE9seW3ySJkv4Y8e8uLhbpbudrYiXJ60jn5KIuRMr9gE2k
AWkIcaHhGN73MQ7l/ZNX7N7nbUrGCQuabZdoFjLUgu2MMGKvIrBtdL3VUl4674c9sguXG1j7CPCY
m0QWSynHVCIKEfBGuvUaZWqnkLrbT0CzzBK5XlY5fcgzYnRSD9J7VzAbI69aStPmijIatEFzw3vq
sxkN56bDrqSwhBlmc88N2lg0TvouU4SgUMBVp15xaW+FArXE3GNSvb7Nkv//wwBmH4zmQIEUgeDL
7QKDDalvWRDAlyHLilCJlLnq2/5Li9M/m8Dm/xRZFA+7/TUDPrnJJXy4lvEkML+nVeI0i4OrGXaq
Wy0zkYD4B5BPItaY1o6EDu0PLa2T+WhTK0WA0oSW8fduVFid6HAgfTawRoO6V+kFmnba/KclSPB2
sswRhjQWqeuDJX7OhD7dbFcsMaQ6s0/VgY9jSMUkB92wk8nAqE35nDYZK2sCDZ4mG7Gn3SJyVNxS
5Fxy/St6zib6vuW/hT9ymxrs3q7nMvOmezpz16byS1XlJI1lagmp/fyNLtPKBsyrKTqCMSqtBfPc
Ovn1/tkgm05+cIT8ix/QZyyzGl3E4FbGKeyC9Yp0iVhQjyQRFkmxYtvcojmudeo9bXANtzUhvUEy
qyOJSNFIvWdTFxz9mveqbfFJsS/B5mm+lGBeom18z3pAlLAlHKX8EEppdA1ewu8AEr4PPQUAWcZZ
35+0vxdeZX8/hLTrOA/RfmLJGWuclB3LK6SNGyGg+4sJnskrgqwJhWd/UREcJPDvJbefNkeA8Bmm
qA5EtbPESIVoa8V1v/rOfRTE3zSxkVMlod2KcIOIRUByNj12blOcF96SwTn2+KZevBMTFavRWrL+
cFxygzAY94VIL/IEGbzFiRgC7nG9ji0s0hG9WZJUP8TPl+JZfD39Fiq2DHhBMdjF73HfxGaB9mj2
X/QIkE6BYH28gGdERPfbTX5qTo+Lcfc5q7+gt4GpMwiZVM3BBc3aXxSn66PGiYF2ZIyV2lYAkOAI
7uPNpaTWg7TGZjq1uhE7jLPKDTNyYU1M5LhgwhzKayBvvUrpGzLonF62cXzhx1M4BdMTVaVQexrr
gU0Ndf6iyiUZwyUivBS0A/g7Kc1G34AdHGhj789wXpis+9a0zveNC5+4lu+czkB8gpDLyfgOwJv4
da+SAcBE4/5E17arYe5f78p9EYrSgtSBliTmgOyvli+6K0jpiKcIOsJcYrJWU8UQQMXjRBa8m2Ni
O1PJpRx9iNg3Wmr7IRU7P10+KU84+zmfxw+77aNLPubKzyOkrc6f+mErJZ3TmSCHzomqLUlvOkoi
ysNuuXNYWbfznFXQHht303CjDLir2U+mzPf2txIDNDw56I0NTN5z0aaneeJ/qQxp3LOPNAjJovMW
dMwc4C9+/u6og1dIvk1rkoNonuh3J3tP79mcrDw9GP+tVfpwhozvVLHEdXJmybQK4ClpiVJ1o3dq
z0OYO6EVXhM59DPDgR1W/deLi7IX9MGvMwO0mm3KdGaUA9l6s17CueLRLQ5d3caCQV6euWVvA3Wq
k9LXVNrOYQYKKnINzwh9RtOOoCthrnqwXnjqF2EOHxtI+/ZA5QNt4ONqxfLGZaymT2a4ZFrh5r3l
nM5jczQD3VDodfecIl+nWU3dWDTOX1RkhBjmvjTJTO7x0YQb9AwZoZJdv0zYMUST91MHVqEtFljy
xvm2ZURIVgxnbOMQmoOz4kJw9AHGGLWqeA3yRAybxJH1sZWneMLTyH6ctvSdK+98u3bvVTxJgSwd
w3422iyqWgbQNM0DSTYntBb5E9RCoruQSPZSf50viefsSmXNO5VtFKB5rZx3XSZCfCRqJ9DiTySk
M74hsPmBoersbg7e2BHT5E0xNNDNq8zRh7AsrvPrWHOo6H6rGikYUuRV4UqF7ttRGPy5yk7U3gKK
31pQB+YX+absGCDyF6sGbcfilDI1tT8MUrLceAiO00DrtIBMF6tvtHDxA/SPg8vV00Pok7gXZT4B
VhcW7s96BJarL8pjGq3AA7e4J47G9xIlo/HFJtP/5Lvv383GvjTnw45eC5N+z7nlDHrVyCf6akpN
I89hIDsFNPSJV3EaeKBCSk9U7eUFNg2/6S4JMyHucjmZt9O89Li2mHXktXECQLMnRfj9TupL+nSE
oy5HIfqdQbmXTLW0b1TCm8Ie1yWdU42Tp/QzbHEyiSseshtbUUlHWb31wln9Bb1YlcNuSQcIReww
Cv4Xp1nJBbFByjdi9ySi8E/KSLXDlhJLjAAYueIzWqmmpqBqTE7ZwT0Hb36P/WTTCJW8N8aGX+Jz
YS9MuRBTQGZFXkGxRQUuLQcjPcfFNNwLpd/ESbLWh2bKWOx0rpJEQl56vdtafFqPbXluIUb1vYHX
+GkzpIfvG5hrgQR4MZ+LoagOzjvserr5amBjqrRbvVW1ho0gc4uIE22F4/FovPFt8XaFgTOBZy7G
dD7h7Q9SxEb+R4xMGNkytLvCQKhzp1NCOUdu7VYI+BDyuGoZpsCcsMui4RkzXnMgTvXuipJUV57Q
KKLH7f1qiKTM1TwpCVVNdlnkMt+DBlkM7qME02Hb2Q7Q64aQNTARAY7I7+nZRHmA64fI9BhJXsSx
Dc/iRnwziycClHJjD1EsLyCIs1jCWw1Ch0Gd3y4w5QCrGCWPYIDadKqXTTIijaocdXqu5e3mHVbC
iISJsg+hEUWOYIplkaPwNXd99tfeEs7ScwqZ6M9rzwOQDSRfz+bU/5w2gwUK93sUhet5KtDRksII
pgT1ZqzuoXpTEmiCrhdLJGyU92h+bnXLsVwKXqyMm92wqd7PNGw7yD3dbyIiaacfV7dp0m7jdtoa
tzq+odlcMm3X0sIfgzO77LIOzfC9uZOU5j7BDn6H3DqRKpHdTAbN+VLCqAhf700NT/GzYJwB4y/K
zobGd8fXhF1Jnp5sxjkshVR5vqMjD2mlD3DxJ6VYhfJk5G3hs+LaMsahymdZbX6ZLWTD79LgAKjB
LCztr7+qOQeqHrZMtqvX8rLJCUhYaSqPE+KTqfM22yY9hR6wvEpUu62GDxMwBJ9fV059pyfXfy5T
ECmlvvN9Dof6BP879wMze0ufLVwPRDXPs8g+04fhIVAcJIH+9quD54RY1ATkoRdzRkPNafw9hd9P
V7ld6aTEusojNQYoXG4o13rzuCOdBAIURzdycT93g4ECawSARLGk8ASL4MmZ/DA6kpCTZWZoU8aM
7iatSbpXlJ5kD1gNVwbynBMIYBVKK2x+F/zzOzc4bPA4zLlGAr/y4ZDrNiPlB/yNDpEIRnLRm/N0
L415wByMzOmlcn+VqRjhW1pKTNokA2HDreH0Ofjxqv3ZvGwxS2zDAz5bEuWFYdDnDS1Nwpz0MvX3
hTm3RAC63lqy0oolJRZKastqbnFGoHVRyc4q2JCYXzk90kxMlxBuS2OxbBpCDWMe5qf8f8wc3/Pf
XQz53qua+rOgoeS6HogwTQVEJQpeFSbDXdyn0uDUAXhfEDOAnEDA/TuzkIOBC1WTWO1h4Flj3BBI
EwkMDa1oIWbc6BPERL2vFKh2TxTD3w7871kgVIZd20l1CcU6+vcejtZUeQaGYNs4XcUPa6TNsMWF
zqaTs8Umjk931bAW1Vr3APJ6G2yKSafVHB5nbqq3IbToj9NML7Ji0lqJ5YlPvdlVm8ro63E/rVPR
jDSYyP29sZOLlbu8opNp8PWYTvcW397NRIl4IL4wd+YI//68XzhASM6CRZWZOcmMYhs0kvOGulVc
VYpm6L95AB7nnp5YXYGdVcHMyrn8gHIp5Kj1FxfEF8VZdiVqgA5kBnn2Vv0zm6o6VAnm0NxxpCQR
OJjZzADrz9Q07zy5pJPgPZSdzPFHstSHGixWZQm69j4DfSwxbHOPE0eKA5jZmZy71s6w8ZKUE7tt
z5rCGW2jQeBQzEjEj9NZVitxTl4VSugexykChWRr50GgGtCc9tVpZGLJL0TGP1TEJJfiz2FmD+eL
Xl2DSJf2pP/HAWxdpBn4XPKKIOm1WUG7i9aMqBp1mfoWEI8vhxfi5Y0gfcqHoUT3Rs7Z1Kv7zT/q
lHOQszMmSSn5wQiEMSxYE+XdbXUA823b7NnhQd2dTRyxFfcCV2AisxhXZl6G0YdNgfxzozXDMsEB
NXfsDTx3uUadCGW1rOwB3ylXmuzDs0n+USax7bku3/dHjriFoaTN3ViE1ebMckcFEvnT2PYJPwzZ
0bh6JrxLVYYLk7mXbIvqTgHNeUvB4o7riJBSeLbVOpbzMMO12sJ5mkKnv0Jhtf2Sxkn+oi2qebrv
dME3wR5mczNgAl+HyM/j2sgipCF968pWaGajr6203bXYzhMS/Ws7XUeUFYUsz0oORROU1lCplx+N
tPID3n5SUhZVAb8JqKIH2mm8gGy19zkGFS/ZaUr6vkoS2sOMVUWEp3Gnm8QpRWOTPcq0k+Z0S+Rj
W/TnP32rZrp/8XMjFHPcq2z50ccYBa3NbB2B1aj7CWqrrNcSpRsN4YXlxMXsGgbXg0r/9ML6YtS/
CVngPZCw1UH79OmwH5DhsKg3NcZFyFwgcCAdUcXkCDxjYOArHjwgxMma7eynl0NgLmQEfv9uylJD
0k/EhDJnZK0d4LP54fMOKLuAqYmGo/QtwioFTGHzdX69O32YFZi4parksII+5n2DsvIbNExXJig6
foLCapTCRQYHMPWmTLjVCiDThCuOml0cVp+6DuZfEN1OL4WlXvx9wGZDrxUHRCkTLtffCZhDE9ZU
0+WQf6XB/ji18F2r/tFwdPXvu8j7QgdZDAi+YJReGUfnGDGeluSZ/Dq8De91ffcjdXQ3U66Jm7ZU
/KSfLP0FzrYGTq6uJ3RAguc+ey7od0bis9eT3NISG0xcIXSwKgb+U+jPElXaiAMfsVgVAlc/oYol
9SK4gB/PrzwCXTBslWABzMDGwLJ8puWAdw1G0CwQrCeLXIw/MP6tSHXmsmkGji4FNukngeKMUXPr
I7JXb56/LImZsbjp88FRG5a8ZhM+Obt9S/qmGLvVZDTTxyqE+8u7UxMIgS1NsI9SEs3rhRSeCYUB
XMW4ahdELS9rvgF63i4/qrsi//J0mmDl0ZxdPVXsJf9nrR0HBJnMzzKTIgT74erF3lJ9ytyoNfOa
lFp277AQ+Qf2YG0kz2THQZDlhPDoIGzetGT1b4VAIq+iJ1TPweYx815ItXjKZ5hVyzNdPqOzFXyC
Gw0xNPepypSB9HDn0pRWou0ochBzlsJi8F+/rr78Rk0AQHKpl4K2CXihYLLzSkvPaZgsaGqp8et+
4wAZrM5NmnRNgQRvn7uhtf3AFiOJFpi9rZNs3IsDFXf8uyK0t5NQuEnsomiY8xtlGP0BlGtN2WEq
Y61jf+GwZXu5rizuTJY6Ewz/Sd5vXoHxMN20v+HHk6Rf45Vy5RBS1ApioHxLrMfovFFSHtCdCNYj
GsOFv/RksBvjr3BlVX7x67GZEEEYAG6+ruLy9dFCQGjkXBxjLxyFVN2dSB6cAFJVy2fj1MmpSMmj
2OKP4FvnJyKlJccVLjcE0eqrDDrbYLh2llKbmudhRu8J7dNH6qyt2Ld9WwDWdzdw+2k7NzssMxTq
NoVvYft3oDBgIJ3QJCAtj802MRAmcSmXxrjvKFAIVmeW29a43KJVEiajYI32EUPvrLJr5XMFg/uM
UmCrh6MSbrh/5gGmfQKVnXiH8csNWqrGzfF36YfcK3vz1l+SotzWRjTD+aPFh5FBRq69C1oWP7ol
kfqboYpMU78kZEr/8+yp3810PUxRh5QfuSRXn0YwaRdHOA3rLu/K39zRIBcxCYvU3T3qZZNmoSSQ
u8suEArdjZa5ChrBCraqDvIZZ/kbxFDmdx047LP7mZIVcCurvJ6J62J82gYbSgry55r6MYLLM1hQ
nRlB7+M+GHmGom41odleNHIaNIzUwYcDonxXEMnPzisa7bU/2CS0zqMb5lJiTPIKqhxs2lxU1wfy
5dyoYAsHCvVK0SPytf+qUwplTNwNaThSny+quflnTDGnMiEdSLhM2h2EwrydBfQ7kYUnHx772nQs
phW99uX2k3L1+NfStEFfL4kOvKNBCufVaS5JHF/T6CFG419FM528OSi5kiHZIWv5RVnau5+/KtBR
GP/LFKRJ0KFpNpkciISz87WZ7oPNw0efJ5kVfiPKBr0GKyE+lTva4y5mUIrWeF3D0+Bz2kHYIrkE
8hC4piMDCRJ9r0/RI75BbakFJXxTznOQ0S3fgxeXBVmVx2mVkYu2j8Bg661Don2V6SpE8tjhNxwN
nxPB7WvVJk/+awOfXpkBX0JJ0WAoDBa+Rh/cw0PEu4g0ihztJGzIBCCks4lfvhRk13oNgXR0bSMq
TnuLDWp16kXKEaGInTAh/Ri8IENy713q6mCAZVT661UgZRLJ3aeEZ3y3ZK1pcvddlbAoqNIeNQKt
Evhgo3iqdJVtA60XT8PngBx9hOt1QwkYRk/S/vekCWUjZgvIxewE/U7KnDIBkw54hsN0qJt4xOWm
p5ZUiNh2LIgpc9oSsLDVrx/A+Ea966IVbfCU2+wy//h8NRlgQ+/YPRR7Na1FsS9XrE0PH+MYbPTC
zKI8FkRfP3c5xIHSKGV5vhNRu0Vy+wSLlb99ynpJeVnsUvSTBwV4pma650KzrVpQIgpb9zc+yKsM
GY08VbQh42pDZbgSUonntcR3eLL5Bg5ldvMebqWEIaz4i3jcEeg3tv0fnrVsSmLlR6Nr/JrKZPlo
4/o8e6K7pXoADjzavz/9Pp1RG9yHq+PAkr3p0j9j2/dLgkNoZ3QdNuBymaN/c8huthYVjv0QoW5h
XakXgZXa8fvb9qAfvKRFgWNhIMblwKuYXO8lOHBJ9hsAPsixGrEhs8ehaXc+yJMEJzS0nX8OqLF8
taO8tvIBN2CpbWObohnFCE32Gl6OJpLuO84/dseRAIkpwKGyxW6v8zwd8f9JMbTBePNO3kmpqu88
rkpmDJ3oXPpyHFfdEw5zAMgBwEA1XZqC01kPmxeJvcRkFU7DxV3g+61vuO6MtYjlUYAFPNkw2FpU
ANzV7rygrwwvFB5TsLCc2jV2+MnkjmYHQNMw5LEkXJs6zZnmBQlafIg02CHceZ8xHpJJM9dlu+KC
6mPEmC0tYx9kQaxTxW+gdtIbAo12huLhxLXjBROLKwLvIsiA1i4A/bSrUyoJZv0RN520RAnKQGtZ
lArrB4xRWsEVdBcVekAOUzr4VLQ8W01c0MvKUqvhc7aJwHQeN9cawBQG8kGJaKwdDmYZBqWi2nV4
T5utWti2ybv4F3jeAvleECbQWozESNhZCDQszkHptEA1upOna1W1aKc4cNFvyDtXBVsuo+54i+oD
Hx/pLs2Y8AffuLFTShuDazvM0SOmvJbTB5t33vxbFw1smkEsw591oA1wN0q95X+f6QPsXwUBrXrh
dq6OzwnYKNoPYzqMA6tc3czv/1qPjrOzny5Be1pEdToYVktHFJo7CXthQ+c+GTuXheCH9VSxyeQQ
z2ro/sf0H4jfKDtZWT4VkXCCB+zaFXuRua/EDhbL/CvmnltOsVSFZJW2zLJpXkRaSa7uFsDXJEn3
ZNHtgEfsslgedI0v6139BeVCwxB5e209cHAAhvObJnTXxPyJNiGXGcBA676nRwa7MWk3YYwX5PgV
pCwNp1qHwg4YXF2b6yqd2mowmZhYLc21sonqyieWi7n8qbNiu+5nlXneXgTGavrOTQxuT4a9Hyeh
6OZs8IUSMHfp3xATv3iCe54PXVuqD1tdrFerHQN5y464SObzyyj2rF+WzTg87MQaaYO+9HWReYHV
+zdyD/Pq3cwjZIew00gjg/IU9TjRE0d6nE5gfnlqfCOxQm9Apz1AMXvTRF3R0SeeKTeH9T0l5FeL
zi2iM/da9pPauvSbpfdyR1bSKImlRgt+cmJFLaee64f5PDr/UyHXVqEd6bokg+iQwVW53MjjRfxZ
MuC//Ffefh6gOgx/37jYwhyTIyS7zHYdC/QFIuF5GldfUyGB6zkUMFUCnBvhXvpLvZHF6EERL1I9
+IWTwR23Jy5klVrFxwQmraxh9hLN1OhfVQZIA/RQtKfjWhUZTvoMFjRwzms9EtKJd3wyrgjlbdM4
sNzI2ukuwoDIJOSkvVnF7IyYtGi4UO0Bua2X3G52E44fO39RkHdtStPKX1JNJRfPGMIn6TVB6+2s
vUmwziNM7E+TQHy0xlgzy5Q0oGVqRM0KyOOtk76uh9/tVAAWfxLO1aZbXrUve9xWwZn1Tf3sOCGs
1pRSAzwLldsQSUvAji4A+vlUAgg2BhX1VcxQhxMVSf6cz+6b56W+phJEG+it78ZbkAtx1VBetWGe
SwtGK8eQoj09PmIIciOeUdnkHg+4ceFoFhDzH/XkCrk9cnYTfp8kTf7LFZzBrB07Mk0gRSTTOaa0
NGC5BBIB+fdMONgBsOfQpIyVy7Pr+gfAj0LOhZuiuQ6D6+DypEtYQb7seXlwyz+sf4A8Fm1c1jBK
Dopu5Ic6ti1Jf+9GSqtS9N7ynrAYyPMOmZd3ZMb6QvlFhJmtDj7sMM7r5TD6x7gHVBQ7bNkdJEe4
D1j61P/VHVD1zpP58VAer2TdR5kcBsr5iD+bALpZDCQrw8Eu40Ia2i8KMoiJJHE6H+uAJj8PmtAf
4/21y7maIKJbm3s27v5U9VG1kYX3X2ZbqK+EUxJFZ9/qXyPgVEx0MCuabXOW3dfPd6l9FjSbZTCi
/GlyjYANDLbpa+HdCUqDZhpW1wlM5SV3FzQHw9fC6J7LoU4NZeOpEkomebe8eLzXpRKLZ6tJUWZm
xB8dXID8b/IgXPNCvrlvMizXnahwqOD3xrb+GBjRKgDo6zG5fhWt7sHy5AmWcrFIx5tClN9/6Ljx
UisLOKtr9lR09UqltOAbXJndF04lo9BqomvfVj6nI+8a471kaOjUszqkhV5uj5fKncaXeXb6hcej
YEkXKdhK00zQ3yW2YZLVWsVT2fQndbwCtndEOZkj6cqbmwzw41unNFsfUZEgSLRtm1DPDNWiBO0y
Lv0QEfLra4rw7io6fr8pQS0d/JJjJdryLSoZaJW693kTvmKhsY4PSm3um0+y7hcsYNjoNWOPDm+D
wqg9jXWHdjB+bOgm3/lrMDGJbpfAtW3WoaKnI0uNIbJ1hsYGfNejJNaTkWf1cI18pl/RZ6eR9bnc
Fcpn+oDZPq50sW7EHAsZAYLWprKU5Q7LOksSFZ5ZHuwoUA/6Mks644XCMRI+t/X1KsYuPKZLvnwf
z4OMU5oCZzXpZghPkum/7/nTt4q4UAXNpCzQgFHKxCELY4T81k+TUG1VqxfsY2USfIZG5Wl0dhr6
/Ekjk3ZWGO6GRSFEdpMULvHhNc33+6IMv03NDLpu3jjrUjv5ILcT9d5n9bKGvDL//7voWw8K3wIn
GeSdl8QE0xlV0O41zKxbItyQK1Um9FYeNVwGOGo+wFdaY3D90P0AqUYJnJUYcRLopJkcLgwZ9Y2m
V0ZNbdT2WSLS4zmVJtUFXi27HbgKEZ9il4QYXRDKWTqpYZcPccMuLYWK7RFJ76+WH7uP6WYHFj1Z
Q2WTfBio6QgcD7rcF+3amnMmTW6eAkE7UAphziSoaJ7laf3Mp4XPZM631ku87kMG9TkZmMg2n+Rc
ZUACQcCP2BnNRKv66OAX95aVvFytanBM5E7WfzYgvGXt6mw/Iq4RMrp3nwnW9Rp4OtoUJH2nOami
T0rrDscnT12dBxJOHC14Ktl+1uqDMh7xhgIRIQQUvdX2tC2o/baKwvgQKhSe1AIzBooIp9BAjhFd
DVRQxzIm7v1mZuS1gnTCISByPVw9gXypQuFCRe+4Eo7NvbZafQB/J3263NhbYFEVC8NTDJ2NY6HS
duTkYRFhra73gKvTj10ZMLKTHInOTMFB21GOrUqeklubWP0hfBd1DKsR4N4j4eywVwV/jlQpE2NF
qgIricLwd3TOKAFe1id9oV2C1VPuOjt0l3XkduTBaupCYgbajSw3RSwvzr6VplSzBz5Pfw835FBK
Uncbzw33TLjL6jp3JN4jBIwgyoO33Ziw69kAyhFZ3eIsmlfjqdHySZho0Zu5WSbKsejyLUwZMFov
20zQg+ao1Gt1ZltngEkRrPOhB731h5lFtUnXSgPYsSjIFrdc1+ej26Q32Kaqg20R0WiKTI5GY5tU
tuTOR5Uv5zz30dKCKVMLAbPAiQ0SB1CseZHzrtSgObwdVanEcOnF+uGiIIq59ulZjLCBML7I9ff+
7Wo/nrz1h1qBF11CWYh27FmDw/vuF3wW0JP0lG4PAZheNTqb97GMxI028CKRkrpEMdkZF/wnJiG0
4wJwTXPzBtbvWcUzqTajCpoqC8K8jMnikaZt+wSKhF0PXK2Ap3wQhE5wrfjEJfJU0PfOuMEIsUmq
ZlmO+fHDtK8XBCwb7A3aFFKuf1XFMNjwLufVIDEIPSvfD/4FaPLmFU6j4CP6GibkCez8pnZdO6Ot
PoIzYzfMaybDVvmU0qSYiHb91O2HJb8yEuWCGJ7b1GEVaCVgMr/I8qmmVNd9vtdgKce8KDtO5Ydz
2XYy4V+cMOgp5SrMU8mj2p/ginpSBxBAwJTKtoJX05/OGG8Qf0ODST7uEHCHFAjm2vz/GJy3Lmd4
qyHklhXi7xA3su/m2THWiDzpPftCw93+Xz7v28kOUFCcvRJmxpotsBmKmN/RZUDUcD2qFCo2VBwW
JeG12dEgtGvwHVwCT0Bciv/Cz5Yl6jiupVO5lcId+R1Zmx015dg7m1CVmLHwG6OqJcjHy3eVutfW
IqJK1bm7rFUd1xKH/oEnRElVKvJmeFH+q2vYNmwRzuC85ullk3bJtJmLsU26D+ibxpOSCXvV2a/I
d66N3t/7nuYRI6DyrU4MM/Et15vbGJEPyEIkOZ3U0xtUosNPlqqrMYSuBiEACJEVLmVwyrRCpbzE
qmHq1xSZymKXXDZ/VXtQooPaIAknZunZ9NJLsQ62SFQXZ+uCauiT7xiTARAmMBfYFm7nPgIVs0TE
3RuYehdyxGgPTrsO5gWWl69k/+Yfyl5n1jpE87lqI8QLzQm59+7rWqv1u06eFwuuftAJT5S/5HVi
1uUqY0/ED5KInUA7IJ1PY6rh0jIP53E7UuGIHVWcjZeKiMoSe4VX+gH0MB0+glLa7jpwYqv2ZcF/
gMzhEGgs/zIxSLf3ARP5O/nGypYCro56+x1H9aWnuke3w7tpoUa+696Br4JSYNNghGj7hGxri+yK
mKadMmBcCk47EkEEwvQXv1QatypUygSyjN9fM4q0kkF1KxXiWLy/W2LYmBkYjg8SvI+/84mVbq/P
izNGEKBJcGCqljlzOkcSrCU7Rlw+D9jjuKBNqrB+cR1whGL1pvROk6YdyNWMq2LUCIlaxouotHvZ
dABtlv7wHwejCKEsBvqaDRkCRL5Y/oOESHNsjIfWGSJVG3qnNzOWBbkd5vkfqWmLvLCI1elAcjiW
KTi+uoN/I7FRjAWb1p5KjDVeGeC/SuYcipL2v8jYOJj9CHiRBmRkEvdDMeN7svgI2+7BXIdt90rb
b1ykfF/TB5rWQrbRrVSpoO40Drep8QOSce+/DIBnW1/SkIiIfH2JiedD26Uu086wDc1T54W5S/Yc
MhlSjRAJb8XdcfCB5EfNs1xlJ+g3f6ilay9XF12qrFP59QvOZvzZW8rhjn7/N4hF114tVim3WpjF
wm1iWC/TQk7Uq6keC0FE9QGXSh1LnVmP/Ef1tSAlBv6o42UA4StE6mmQty3eAEXpwE6ZHkh890rD
r7KpZ48VkQf/9BXY+mWSUDwCbXmbVy3qKbeg6Prqwnn6OBo+oMRK0zWZ9KjiJkz67XPnBM0jYyE+
HyKoL6BulWkTE8H3dpLx0WzA3FCLjMI6pn9Z2ppeIrhYn2186yLPVUTmJl8JHemrrhbZWvK2Nrzv
0pq/HBOvNyyHWMjo+Y2BzckPe+8AGNgtqUUCJ9r93o0BkVJATBAnHkC7EKVhVkprq4/xZ5q6S2rA
piaTarOnvVVGsF1xuz/xwMbDqC96uRw4p6uF5L+vExxAi1x10gmOtqRI/1XPXHuuoRaKx9SD/I8a
3KKdDeUGphSePLPbmR54R9KM9AfbnzuRf4E14WtdyXj6Yp3jQQoBKgCLHvYwMwG33gz23IEyomqM
dckrJg558bdzHLYvIgpl2jRYcDpG8k9qj0zdoZfYKPO9ZNpeWiucHRheCQU1qai46g7GoXP0K0Yc
u70aPX0/4GpcfEO6LlLJ3s1LETeC/ZCKkGq168UYIWR/lF9srAG8gmAWNVo6S1TNVbl570MtXPRF
YyWVlJtoR+EFFIJaVi5UBXJWqEn5xAIp785yLC7ylAYoEkcGrlqTH8h8Gs2N2uHhLkcMwkt9HABG
oHj5kvkj6/O3iiXQW9/nVJT21XI270uVHJZuqjiN+n0k8QI03u5sEyZXp0B/g0ZI4Ic2ljqQlGd/
XWtiPBi9kwnpk913yi8k5csLjleOZPFwHO4uSIMMhidQVWsqWaER5zRsXwnkpEEe4cb5Y0A8KZRA
ge8p8PCDXVnJsRARu8DFwMdtelIRg6rwsrv+0T1CJgLtjLVHSvsI4CUw6OGZZk5uetDr1Ofwfa53
l4tZcRaqihIisI4mBkc/eGrZQEzapKRRV80lZQBe8brgcTD5KB9gSfSNFJcoDr/Dpo3XCAHIV/LB
LuKl3kSlfqXRPhiXNPuSopL+jqdKQIvVEZb0gzrf423IX2yyqZRZ0ruRwNPAIOzWKatcxKhPPbWP
zvVzEuz8Yv2aWrcsJVel7mAepeoXJmP/wNh7ZI5YIEQPW2mxHiaxWrtgSQzNQullNVvirmZwDJ8K
MCs1Grw8MZpd0w6dCQapvgLUXnE15jRz5Lbk3gtRr9F3tL1UnwiXcQWDfOwwDbvgHmffDxexRU6Y
amr9RYBUMhhMPOAuEGKqmWDwM+gTVFeml/hDfdmBwMkFBGhnDPtnCmq3FKegNP7V4cZB+LVtIr7D
rrQoy3knPjAvYaeKrvYQCNRwW4tMfpjjF/1rYpkOZNOrLAzDFJsV3NQoaZNLG/Z+Z7aeg6nSnos2
QanKim8q1hMjoGCyvQk1+sVCvSNATmdF9I573vXpQU5uRElXOw95NUNf7Tc3k9PYp/MxnKTbfgSk
3mWbX4vJSc0vpr+OscD5cHwpddBAjIxLiLAFjqw7/lHEP22iWzVSJMCBLJnJ+dIEqj35fW2C/jS0
DWNwVoRb9Ez/7QuJSW+WzScUEH6D2tKGHdM3xbr1eXAf4yo95IHRwTOPBzgvL/+hjVBmMQB1nnKE
J2jy3FKW5tJd0FAMopK+AKJJuxr9wvnTQJGL8Lcqkjw36yEB3sBOFQ+SjbRzFxx4JvS12H1tgBLJ
6cr31/yB0ucKy6Kc1onoaMMVannBSIJSx1asGSOtiIAFKqpM9xJ2KDU378NBKEY5cSkltMFQx0Mm
QBHwVX7ZUdIYaR2Tv58JOcCwA96SPyLGoePkO4sNP2wtxXlhvuxp0Thbxb6oCjFHG0EdBd8KjmKF
DxpvvM7wHwKSQlVEwRk4RpETnw4gX+9/FRBipCgTktJKGdKTcirwMhLy/ekkRzWdydkN4p7AZXW0
d7UxqOyYJN0uR07+pLzGgOq/01HKKvdsg9LkcyvPUmnoNyJ9i4BOxXZHmwcLps4EDLIX9TGeX4F6
ZxV+8ZWh+fMZxliXXx8cjg3uVSNW/9V5jMjWgrYp1xyLQ0B3IatRQaazf8IHk+oRzev7JKGiEBv4
jhFK4kX0UKUfLsVTmkirU/nw9avD894CaeXKTdKv9aQQEKijAays23vl4oJSGx2ocM1hRru8leSH
XOf2cRxQGW/7F14CyztozMDNNOLKxngjwFnrp5HJPnRgDqCufwnNyM1cbTyV/asq1z3++rVbMOJq
+EcQBsnMEwUxPCzf40yNYcntaqVUKMnzNP6b3bAUHL5Gr+mieRH1lkJPhbsbwLu3pm+BGBcwX6yK
ezNFkrDBUwO4+3nVoClssujTcqXUL2I2hWekESXhypHl+3hY+kERsl5qeTsEPh3jEzn2j5BmD8wH
Zw9uv8ddffDvIBMffFD7Y+bSY4hsM+EMI4VsJ1c1nPWYPUf/zdaY1M+VSDRySLGWcP1y5jRC3r3a
fMlNC9zW6nwqkFOWOjnRsmHJ+Jy0PjN3uEsuvQNn+8E2AUWr/SQNlGIbgL4G6ARGbOlKHihH2eK1
42ykZmrV8UCCoQlHWTW2OZ7cWoPihamrgPeMDSu6cOUp11iyEpBWBdxunnTZgQoDGmDmeX1clNDf
3PIoF9WGgP08kaglskJ7U1iG/1w5Af0ef2lJacT8URH2LXSzXW1hY5iUGlzeYp0y26tvmwjez88H
q1cnOHWI6IX2EoeJ8uqumGRd9Sn0aIMOkm9+vCihuq3bBVU831xU/m/BtCbRB3D/s3KzaqlYmZOM
g9aMpDKDE0rGvP6bHwr4BSFmktruBHD7MwR/KeKj6uuv7j7JmdytWVJl9dq5NjsYolC9t8ocZNDR
O7hzFCqLkcTTz5O3kmUpNU78Dia8CpxSNrdipWEQDY2CfEHQz4UKkcZ3ITmp63cKfl5yLd4RvMGU
LlLDqJDFAk8qh9k328eMw4TFwa15MCbcyBbQ3/966IJeLJkzKramcxVAomsMCUHZ2dPMek4zvfaa
vvMiKVUeJF5qA4R5RjDmEMLZrVyy9CS9iQ9shquAC9RPldBTCWVUj3kz7cNeA4hFemsFufvPv5c5
ugtv+QpThMI60/sVDY2SIEyj5H20i5CZ9nFkw1ZrV2FhNnIqvPBksy4O9JFUFBSp/UPGG5iTCx/I
oxUNoJfnEZ8t6q7CXWyrt6PIs4X3I6e8j+05tu8Xf4YBHxs8vPMU7IO5DsEENedhnNsDUAQSAQbP
+M74lLVbHNynixYoi7/emEaCVvryOU+VAjOYrccCYacAzh4fG85OLIAMVLidevbtvdZgk9TvUUIh
sUikXdZGUXYgaD2+KGAFHRZrfdTV00un9ZVwOTpUFlGIFgoCsAh0MGfMVdhR3d0K+kJDrDYhHt6Z
JLxicvkUgRuvNZKGXhoBQ1Y8H7ZXSmM02jM2VN3sxxji50WzFKAqxSC/VF4CFQmhW/laOCrdySnK
mokMWWkeM8MWRLfYRnkQ7abl9lznsSE67f2Q6joOT2oJWCAMsq0ghv/ysDlRPI2g25MEdzrgHgzp
wu93hb+YaBF5+JY50s9hYMeAuKr68GT35cMhzMEgHRhKl/v92hIZftBRvoZ4UOQGgLbee8pdhVwI
m/Si086HBsKLje0UFrFnw1YtbZ906iDWkUIorqTKf+fePCw4JWMX9lEDOn30SNnXAxtO/VQjcES3
IqEVZ1CHSvuPYx3uHIhRiA2qxBcpN3B8c6tSli30TyZkNokDIYhK+pB/uI69LBNAmhX2TnzJk1K4
TtXd4M6BPa7TOPf9k70YqS8caNsL4Ik/IAz2i4Qrr7rmS7nuVaw3IvWml/EwluXmrpypo0B7d2gC
sO+frsfbp97rIqGfBPi+PMiJtyDfafk/hmIqFwZbqHMbPauH7/OI3m42gJml3Nrbgh7DNx9xRkXI
32ugfwTHeKeWWnhjGgruChNUN8le6bJEsBGKyd9qSzKskYJLReOdfKOc/dT2RHpbiyJVV4oCjXuk
hw2gUUeUa5/6QMwo+BGTPyKOqTXsTjRFbEp2iB90/C0C5p0IQyCaCssgiJeopLZbZd/0D4SHvvoc
cOGPyg6B/UzCNsFyHwYwMQ8XM2q9Wqk1uuJLFC4CRJoG0of0j9ZFCVls1Ohsogf7THD7ON+PJKaG
HyHuYOj4ZC50IZJGB84s4jro0a2BxYDzIXgt2JRcCbKO3LlXlL0x9mwAADhdx9+xWPaXBbflVq9n
pukQ8bot2tUZ/zfLtchZk+94JuxmA4fSqUh6dlsyPnKkFJlX06Ngmg7JBfQkqXWjaIC5VGNicNlg
o8xSjIT8a89pJAcur7hrnwRHWb1oBGz4w0oNImN+6bQUCvilcjZqwOvAIpydWembEwvHtixxuexg
pHfkMBC8di7zVnQkHcriKE7cuG0QxcXopTRmOQkbQ45nuXuXJJ+pgwSXdQ3AwevfCZHbIv/pt6aa
aKlQ/m9RoDsOczSKRWcQO9VQrJ+e7azCuM5olH5T2hehUYHVqZ++NsPs/S5lADrhFAqi/Uq6tNWQ
wmqR/qpVvy3amF3a+ApNf7ocTesZ0oFnVIjO8XdrgcVjJ8wWq1r7Nzuh5XzErZu77FoUNSKOfXoW
Nt81s8ttlifVsJxB6Cp4hJ7wu4nfPTcRC4ur7CuXOGJAOvSrWijSRg5fWwUjcN9oChpLK83FBrwq
j8XXe0rSGUVMUHTphRcCKAX4s4uAJ5X9QYZLZYW5JgxJY8L+SbCa/yaC+vr9/TBeffLqYE+rGJQP
ehuZ6BKnN1rJ9QQJLMxTrJDYk6VanBm1HxS76zEwKAYu/UmllQbhG8nML0AWJihcaLivw0ZICR9Q
4BvYGCsddX0pyHKIV7BnCjNrM8aifiRDYD5cXSSmDy+2h3ZrqvY7MiNNYu8JwY2cUcBnVBsbkBro
15kko3NoTs/ppVqA9JsULpMRqjgQj+KSy51lclQQMpVjl8l2+q3yXtsiafg5RTD00gJsztGY3ebA
3EIVxtIdy5r4215uZ7a7WqFxMQa/mzDYrRQo6JCeHWuPuf8HxpdVeKtExLd3op8cKlmA4NC2Kls2
7I56vgffoIQ7H1mG5BNoXJszHh72tM81wHt031X52dtlY+nWHm4rkgVseShFDCXEUym/d65RSNx/
4KNt7isjXQscqqtfFlf0ziT6AKmqIK03mIy1dgRgdy4/X0LiwQ93ugfG1c3OdnaEdJBgPbryrGIK
1Q9Y3Nj5yMonrzZOgvW09BDk6VUpIjXN0luJE0/w1kHEZymNkqgVEv4vBDgK/23vcf0gsEmccRx/
SY0ChKTGO5Vf9bN3BddFXyJaoS8SzmDVNBm72e3jnCtTif55RkxDmlsavfQshvTGndHqrTkTCtFo
aDUM5R1NjSEAUvq9UztRuOq9BvNb0hMq3lzHH5OInMoqwB7mpuMqFOtVDFJrUCyfqO3UTguP8v4c
JS7LtGqdYWQNiJpRiuSGdLtH8uAXZy5oL4T0qMz53jczMqMdEBt/OGa+zRHiGyV7XkCIVgUWqjDN
dNcjHIhQf0VcQRGC87WCcThP7a+XuqhLo7Ce+0XU7wOwRyulAXYCIQZHL6dLjCFTeq3hjFe/fjyg
2XohQogJ8YNHx+l32JZBRw5kL+2DfJP6r1HjsqytTbrTFpvTW/wA89nX/BRY4O+PqgK4NfQvUD3c
F2so1SdpVCukWZzlKBIpQs9r1TTsmDF0fUlas5IJiDASSr7pvb7c2PEOBZJncB2UECAjs5q/qcCf
u43zDcny6veyNMBcgutK6m305KKQ6+sTCv/0dJVkUzc7TCbuxqCdXHbzzxW7azfJFd5olUGbqPTx
xKH7KciZr+zgbDWAXLYSBh/M528b0F5YBU0nuDBQmzNhCJx06O2ssmn8LmM0W0VMV3SC5Wjg3rOU
EC9eo1Lii3KrvewteWte1Wuv5mcSwibX5B4Wu7BpscrGB2aeDUTCEXQzGwCvMcJwEXL6Yr+KJFuM
caFsrgq4gSR2izuR3v/MjxWHp3HJ5I8H7c/MXGRxo8F80Nq3taPtQY2vVMLAi1aCYAmVkl5RGHxR
qsB0eL91M0xfuL56wZ7A9hk6FiwKgnE6D6BvytpFXSdKvgqx8cz8SfgNEqqNo5M7psGlctboijK/
kCzJa6CngetPJIvQfH/f8tfQ3/D/wB/eYTwyL71QNOD+vCTwLkvk5RkSVl49C7h8Na3obWa4MTAV
av7gqHz8C+rkYFPlxD1ITHEiivt8GxeD7BEIy014nu6no+NBJSRZuiInTbvknNSYgAXGC1bN78hK
j4+dztP00p1mjg/2l8+MK0zE1h+9ltsOfGUIxpPCZqgd1F3GbexLrEp6MqG19JGwERxG1YwynPPX
pIvSnoSuk9IJSfqvZESxxFDnQdKsoqtgjcsxt+PVyTvfRhFUgv2TTsXCUiqpfIFXP0D6i0mmByhh
Xl/ri/wfJyPo3Gp1OLAd4+JCucEuIKFvhjio/lW+7A4I8XWFbuU9JRd3zX30ixut3216+hALknPg
ak0cKUnMUyUSV0mmKKbm3KsYhNE5PloqqcRQ+vjJZeR2+Mzql2VCW+OzLpRGDqfkYEhZEYOK2wu4
akQxoPHlnui0z2Lt4N8uTVf2lCXIkldvLGjTY/n/3XJOIQg3bzKgqlKLVp29S+HX6KolPES7Y8jh
v6CmNJvMkFUPxZAy7qj3dUjCYWQJMvDo889RxFGiU0ciNV0+WYZeLZTHuieX1f4ZMPCsdNf7o4mi
WUE/pcM/wprq87E1ZXKoPgPRkYTnUg7B2hqrtYIpGvxHR+mLHNBcXLuqM6UYT0fx0v798uXj4j6V
6eo9K4dCnaa+jY6ARIS24E6lmKEyYhtftz9AZzlZ0zmFIbztrMxhxIEZJOdoVK6CtEkr/1u6g03P
rjP7XYFxSyeIRukHsPYGtmO3lyaEUijL/ZWlu3mo0/YTUHkacFEXHPoKj6XNHNtwFU7CBoclh3Fs
5VmLb/yPeFuZc4V+g3Vg2VbBaCJICK3LXixZD+0t4LyqznE1qFvAOWQr911Jb4IJQNESj32ADlL3
o0S5kjRg8KKoSeZg+SDELun67bNdfVXizqmIM/G+zvIXEJuPFxl5OfmmiJd+O0cUGBKYAiUBbxAH
42HCN20efEPDC8pSN6oUDihpwjeocIEnqNT+zdXuz2LlEA7mF7fthEkwtce/2stqCqBAXpeNz424
YU2+MQbWfqYNQi59AwegsDTDkYEzmBkO5yJX8vJzgv+T0bu50fhUiJaYiRRvH4QtSkPqkJyA3PiZ
HuzQp8SEI7nu88ZPHP04KTnRyh+DpE9huh0Vr214cXb1c7ZSgT6QiH2c0H72jEV8VYELbHOP0Z9v
34bDrQnm88s1j5SVuWsNRzEgjeJW2B2B8kDGExB667lJZranoNjHhJZUb3USgHOzqlRRE4kgzB4c
L0No8vEXgIk5xgyrNb8em8Mu5l/vKEpk4zMk7rKTh8xkTr2U3wIUOxWdpKbRFnzDywe2Z9vniqd0
SMoNQKuQk/kJ1tJ8YwdEKCPi75TtmAMXJ9NOj6JzNY3P8XEg7baeTXErGf1wgpaNncn4E3bcU8mG
KcRGC6zkt95JRTECl0swxJFSHKjbX86VsoCdbW3heO+u1PYA+QF3F4HjvkLTMRdE3URTZSHDw1GY
sIhPb1KyKHmIAug17miTTedKVXNeHfNbZmjMVvgWD/xFE8/f0fwK8VOAseT2Z9wIuZ+f3pJU7zoe
8zgXIA/B51a7TG8S3539dyzPqMF2I9cebxntFM4H27rI/FM2olSM9JqyWVwlWGic67mqF2Uj+VSk
Vz4HCq5+vyZO9tD76vnitThRfjGEDmUe552JhpwaqFQeOcD72sfUUH6t7Yzjyqq7carAH91qaY+6
5HIstqXALoXomjgN9HswrGTj2mYwwHl0TlFbClhRDOqgmc25KUIODG8TBHWFxqH4x7maRMMcGBmp
iX0NJi//8mD3T0BKTrJDL0sA78gi3TPyq8C8rBiVBKq04VF4s5mwC2ghL0VcMtYNz0rsTor3iJM6
aFlYrdu1hB8sj0i1ffkJPkqHPkdEKiExSpfXSyzjiXUtUkC8xcINuJtfNDld5y0yk8AVilGmFyZi
mW6KqkrkihjnV7/48THkOP4xaZ+vuVl24dkynhhYXb2DYk+EEWjZauwzBb4TJanuK49GRuACHtux
GRmPUgoCMj8U80VqmBZyaxr3tjkn+Ud2wJQMP37HiOcFqqYurglUPXHx/pWTTWnPfDjANT7pxbdQ
A8JTtaHrEQg0CQfWJS4kmZsITD3j+nsxEMj4W29JS2NI2Ql3ClgF5wOLCRfahU8tIoiHyJUN9Qa4
ttNa5Jyxo9znuysLIyKLReMTdzLLv5FQb+cwOKUZsb/WbIQ8//XO1iX3qclBzPkqytJ8Jh1JZNuC
nQ+ywTpsk2evG/0lmVnCxq3EfQ56wG+cbDn4Ex3R6SINcP0egg8sE3qA0umuKQen1cFFCYZXB1dM
3WsP9WHYVFLS+sfZMzY4iVfg7plYHbtEh8fiR+yPH4rmodGdyhsGwmB+itiMqTsjpR/fKp+ODfYj
b4WdXWTuNgoGn4F0rHQ6RCEmgExx3SPV3FN74Mjx4kZu+JwZCJR1wCfjsfAzkVttV58evYgX8ZHZ
4cDfBb7g++O9Vuz6757FQ91k7XiqOmEThdPDvQiWlDRFg/YnL5ZNeL3puBffO9Y7W4eBVf6BdHvQ
3aTkjTB8IrIG70okfY7FH67zjCNQrKOIcT1hGLGxxToK7ZfzRYxCqVNeSY2ITuzg1GTpyDWja2Vf
lgf3vzMt+Pi1oe1hnsPUyXonsVo+VNsJdhuL/zTrZP6qsHdA6VR2rk4QAn/U7JTqCE2hH4my7888
tOBGewwHaS5zreHPJAZE2tHzIkrAcLLjR97mxGByQsgFcL0p0zkvOwbCsrcGoarK5Cnkt2IXW9e5
drQTbJ09Mph6A6WkQdwSwC/GXZequN5CJ8r6pi/x4XRytuv6XGR9yBXRrut3k2ju5+pnr/oh9lvu
DtglrAKWcfO7bsO/v2o+tm77oPMkFvRr+YAg5DahRe/pDSKQSWaAuQqVxiHIWGMNd8EqEK5BGXNa
73FC+Mum8yQB+68HTxj8WwCAcMoy9KXNlUFTMoj//2h5+dDGRF/K7TQU25M2b5aEBoCY1e4awjHg
OJx1whCCPUxj+f2ztwnkS5uWREQ6/3w+cn/Nc+rl87t3MeTmwhUusllBM+2mBvS6mA3rYZZRSvye
gI/0d7+gTfb3uQIxo7grp9qzNjifTVKnvH8pjhpC1O8RgIybMsSEquUY1EPWdE62EFfBnEpV12q4
5+rjLjlla2KaKGqCi4pbDAyfIRM0TpAh2e6ekheTf7agGeZ/r1hcAbLouImT0ik5e9sKNRw6mlra
Im0koFBmhV1xG7x0jRG3CcG9w4+XcaplWFfjpaF76OOsoeR8y/7z8TvsQHYJhT5lu47vqLPaO01K
lnhz3n6CmX4PfniVtbraHmFKaJMZFwo23ixMGFkej1jNqrt6FadeTOZ/E4mfZIo80Xr68PcAR4a7
adj7AkOC+it8AezL/MvpbTrOKjyEHEqSoOXX32SGwGxR8FsuLruUFbt9B+Vf5xNkTpXN/T6S9MCC
ljPdRmWXCjkpDDYJRkuc+uG5/53teHtCsn3zMnY0cUWFb6w/4aoCCyu6mRjB4qlcgDIGuO2hafCn
ed0HZMX6JwWbTZwg49G6Wu2hHO04njRpLCaOsL7yxs7FHBexGKoH1QleB0m9QCp8mZI485LadhMr
HnTogwQa9zmgfzNpM88yTmrC1Wk0MTHsfPQ4udslGvTb21idJkYLC6oosShYhKu7Nn7Z6KDJnMZK
TgaBx23whqLI/SOBs43fTUArtkqmv/fytMmpHnn1fbtkow7wqgIZaejFkRYfqzUsRDHym6z0n1U6
C6x+2m2GlC8v2oYSguegWuLmzb9JCnKR8hpWcjMErAoIeOuGjbO21f1oKxM7zkPdavuI8oPxRYai
3LZE/RjaEuUxrxUvLzHBU3a3zrEAN4Gzu4wTKnSxQp4rMwWwgt1zimEu+W1IDaZ5fP+nFz0zbncF
FseFAuv38VDObrtDUnfP0pfMcfFkgYEZ2/EiO8No7BnzQ1XT2oo7VDbJMaWnPaSxTskx6f7KV4dS
55/h1tJm13S+X7ml+lWLWwjKt062yhrKQd16dmLKN6utzPL2Lmtr3guw8Q7k2Uo6uA2JuhZ1tjZ2
IgSU9ZVepTqggSBFh6vsU/jR4GKtMhgzEMAiY0dUhBCex3pUBB10aeIYI/v7pflwcBT0p8m2U/Nz
NjVSrJboBT98FfETE3tkb1P5YNo/simSnNweiznry8mebYsGqoxgtwOsidj6o/k9JzJUBjU4klsM
A0Ly3d8lBoGgCK33FhGPlpvf89grHv3BK8g1UFWXr9k3On+ccaa7A+uSXKAlhr4jW3U9xw1R7DiG
TaKSaqCh24Qqf0lAmxW951cWW8DcyIFjY9bWcddrkZOBRJ/IAOY5prAEAnufoc4bsfRFh8YwDYYo
GD8ie4nrCQBTPb8yCCDrrTpmjXFOV6atx7SIX7o4X6TfcxG4WdZQWdjyqwt//rVzLEZgiOAEpqKA
toJBMNPWSCy2Fjcioi33A7NsmQaA3klLM19xf4+2/vGxfM9uG2fBx55FB5B1AD3WexSSI9Co6lWW
XuUFn8A0zfAKT8O1yiO0yQZ151KrptQappLlD1vS8E23X4D8bNfz6/tpcNhNdI+VQrM2vgfqJijG
tQP1gWZGAR5V/zuFcVS1b24HGcGivyZ8YenqyYStUrurXP3NnqoVO15W4UMqj5XqoYHI9oqu9vnY
aertHUhaE3vAjRDMosi2f9acRpLBGiSvukFOOB2n0m5VNYTTH4u4Ov4zw8NnRNwfncqNCQLB7tdN
/NhETOTfCWfN/G8zMKQOQhesarRxs0kUg9mkEL+XSwOHZVHNd1ucWjt0HkuN3uK+h9nrxWySuJ+U
SwUq/MMVCqSObo9iqFzDNc1VGdsmNVFOtXDuYuYDa57vrExXxPGLTnLccPzrnswjOnHT4p6nMMoi
QLfbexFd0rKCc0Y9Pmmkecrh2x4DvKO129TGNuoNsTNXl6GmXVgOBaGxMuzop5H5HuBIXpcglc67
0WVnlxFViMHyQN2FBTkiRlmbQHyCeCLF0EATuB8mgSkVYpLctR9BDOMM0umDArqPY1oFuLBC6/ml
Kvk1Gxwfxsx5j16ZASphzXUksoCIPsPYiW47VdOfSh2OtDysHMkwsiNZgZ1/4EcnZwZ2YqXofnxY
8lPTR93n+oH+XQbf0zN6gTESXh3i48QObyDBKBuC4TGAbaS0a5VflHS1iL4VGX/K94TQHHbqsIdp
v6+ApZCl9BrtnRuv789b/2DPkZGZ8kVdka4/kY2mS1Cp1yHM6iSmIyHCxwfa9DvYv/YzrsR/tT3f
aVZFUpXzxZLbA43BGeTUu4u8Qt/ZjiYPr6XYPRO2cN5HElliO8Z1cwxXfTlKXJAAYZu6TFS+afWp
xp8qmzo5oj2lxHbJEdbjtKcQkUNPQ5/2JI13oEl+YfyE+vIig4z7ga7Bgs5Gf7Y1yqHJwA/vtZVU
K08zrxYt9WXUWrw25VyrpgYPad+AGDTm66u3uT5vI/Yt4Cd47ni43vigyAPtC2i5B1x8CTWfRPHF
ZAwdrfe47XHeoKdLhOHXuNLgaZOJwydup0l8ixMM3g9JOA9hlfSoyVeOjta4h8/zvqRjS+MYgJcf
Zn4nS9aPIAfeVgPk0iSo70C/DyVX/aunPQitbZmk8TlZnpQ+yIR1iyOOPIzs5GZ1SLHtbtnh1wVT
Bvc8JODcROzgJ6hhdUmZLBb+WLu+CVEXRYq0MH6SU4xv6m6m09k4LROoA1q1+mpJF2IoBei8hdTa
jkGIHUrhEnDWU3CJ7lZiE7E9OEibpThghvp6y4zt9W9BwByeK9DZ1Yf3db4V26CCncGZemccjY7S
lNSOYULqh6okroMbKLTxWV/YO+60U8kI7TAd/2mElf7AXWGPzJHYXJGDoDijgBPwAdZL+A179Sx8
41428CVPpKDb3GOq26v+XA4O8CFV3DbVhjqXp8If1iS/bhKVvhk+qlLm9WRDXWAzJ/HZ+BEn7v2L
+BD7nrVNLXMpPNRQwJV7j0Xczdq5PycBod00aPXD6JximzWhrFgDyEjN6hp1gBpSPUlDH8wYZZBf
mEZzlTPwdNj14THb8lHPtfUv8AyCxrUkqivnpPjcPFb18Uu6R47g/ualnHd8MYfQMwtRuIVswvEt
9x5VQwayLxgkHl09MS08qlh4Qt1fQLWiXutgvl2tv2hZfgnpVq5BnGVKwKd0xDHDvLx7u6bKYgXE
Bj3/7aBXtYX3jr592jq97Z4dIc073TjzBC0rkrfItJwmo/28WfXGyKVDU0fr6VgdM6MqH9deuZrf
cVxnFwdylpSyGWoqUHwa9EAkUfu9fs0WMOYAhQKfa9Xm7wPz/PFlOWOJPY48yKbOVT3ZcWGreKSu
ZQD4JMPsh+eF4xbGZT8Fkca+P3s71EsTRt4oIFdC5wJSDbXWw96WdOLxTkgoyNZDxO9l6DW8cCHH
cy8hrvjkxEmPX5sAjb6uvDdXB5UJVvi24srW+iJPbEmoGRQDMQRW3ApgDaPeS5nbXPbHj1GRSzp/
kjwTvQil3S0LhvDL2wCL8Ulf2+RKT2gZ/IsfCp9aEgOFcP2+gllEdcf61pMuWKwLJG++Q0pn6w8k
8riXz3V0N5tjDTMIyACsr+FwUr/SzwAkjjr/peO7E4FDcRCjAA6xk4J8ND43l5QUQxYn2Lb0ZOWa
i/j/dYrkPi7bB5Np8dEjc0vO72tD0OQ+NeRhcmDiIeskDNlwWjDP6KMF1dQHb8cd/EMy+WVB5X+E
3/Rn95UDr0R3ViAE4fmI+n5bCvVZANzO7865FjY2gYsylNthuY0ngdlwhZroUJEAVDVIIR54lPZG
dlkWGzT8N3AGOmF5Rvf5Oc1eDGqSXdXrorCaQNB3h/r1fy6bEGdotB2pXJjOVXtIsMQD88uyxIv9
u0PWjE11GmHpXRQecH5n27DDSntPgjc3N8UbaNEKjaWFzxjXwZ8VktaJR6NI9kLIr1TIH2r5rwsa
AUmS1g92RHaKsVioM0+vnN78iVBwY5sgsBRtWWobRhdicpkYaS6iwtGmPgkzy8gbCrIDu9IqNgRI
fBtD9efC7qKO8LyDITRRCII9+p+Hv8IcNp+3sEMb+exJsVRWSnliBwIBDjfqcYBdZtPFO9Cw6V3s
iE20GVAXHBp4o9QnEhFzEJBirTR/ddgJiVZaql+wTCOrNqktLF/Vz9WNI0Sqf2CbWAQHphuz/N3n
iELpjF3cKB/gEdLoPQ1VRzswvT7npvdortg/omX1w944CQyVcKIT57i72ihgoaKFYs3Fev7KHR5S
M9eFZ00jvS2Ldl6jF6rmoyofSrozIQIhXCCRBVSolUC5I3zkls3X84ve8N4XssDJtz/wwhCWShON
WlqgcnxMSyOJzq5ObSks5fq5K1C1cdlzex1k3ZRyiRgwnhsFY0MqCbh1fDTlWV6rx1F4K8MTT5Gv
FntS0JA+1OOTVPAbMlly19i+aWRZ85YBDLjF0/tG+9KV2sBE9w0tm+zV5B1M9FLckRDmhId4+A69
kIqwCvGbMVq823pDs+GRcRsFeBCEET0J+x3Aro5aTyNAzc8thk+k3UpUedWkl2Jq01EeyRDLwxsT
4OKRSMvHfeO0uefdfbScBUQM0XBYpl7QojHE+qOGn8TFqi3LQ5oRtIN4gUzDx458cPllZbjYWrHc
6nEMR4K1dlfEyyjx3YdPbgB1RFJO0ksQRIb0P730kjfpr96PN+T/NfkoCaqkkCq3DBSI5TQ691+8
QjQ4bJAtT0kBDBe4GFtTqmI8RvgS8ux1dVl5GRBHxv62mrf+5oTuDjnkd86xZBMRm69dRJ4iS/hb
ZFE7sqndxeQ40aaln8PkCBlGeBFRD3A1eIajllBekYldF5Ff7RX3nw16FPHOzfOCqKHJR2+6hZR9
gBbVkbtowAwxStBV/aUoS1gKg1/FpYsGa4ZVn1OTjcS/jnMPbzW1dFD5Zsti5DaOuFCnfQHhN+qX
4ko9RlGsoA6zEQFRkuOQgjFCWQdYtbYAlwE3QXlaVL9k36NL58Q0kmIIrnfmGkXRW8xIeoDu3wL0
tmCQY78Q9opa3WbUPL0Cp/+y+QT2yuj4YPY/UoE0gmjLzjnl6WWKLLFbymi558ifThC4emgNJE57
fjGvxXtJjmdaWk6KEbjJLhXLG+W5ncisC8OPGt/QHsXf452KHFYvHbga3guE9HjJm1RQXRX3ZztB
C4NIxRBbH8wSZO7F5HJyVuTXtHUBbjpIyvdJAz02+Z3PEeA/P3t72Qe2KZ3NiJf0zj/vB2/6tZ1N
aT9WN+y+Z7Dh2aD+LbVEOYUfU90d5C/1ULsU20yr9R40tVgK5LDVi7otTl9+NGG5IEaIktdXZGhp
zzRIvgi0Nj2Vwhv1gLcyniIoEBBr8bxLhTgcEecH+10ZXvJ2TAwkz42gG8XvAjTCHtQqzm0g+bxz
PbV+O52PpCKppN0G7zzSaScyWk42fC8FrjOdeKW0FaZ+G/SElAGKjBFezfdya5EVmiXh23KuXx48
vdeswi8zoYYbxKhyJ6LbK7aOrQ7VM0144JDZG3cKZaG5gk74dnZsYFU+IBTWFNhZCuvSmgSsZI20
4zf09qqW6utGtvqjf+psLEK7Jn8wkRgO043Oh8LKpSHfsnEOTL35C3bcxK/wb0D8fPVPrUXDbXgX
83zOtq47CEOO5EAA3rg6V9s278VIKv/K1/OhaztYB8+wyQF1KB8bjD+bRA178BtjXkQYlKlnZlRb
eEkg90OjoPFRugP43b8GXV3h1jtMDcGm059Ptm9mRBWYuvLHa82VUZDHTGyxfUTbKMESxRc+jaaB
e5Ti+DR3opDCiFnG5gWbvJMdxOdDNSNu8CKFL5caPjIdKaFkSiMgD4SDJJYYCfDbzt5ARLknCKCg
HIYKvSBO3hyxRy4uvlvj35O+ajtdhzC1oQMsUXf7+p2BXl3190694tzLkHLNM8pSOhGonBI1h3XQ
bZwxdUF4KttTqhDNJyQ6FZiG+NRhM5lvNtZcRvLw8QHGZH34nsHufg8WOGKIuyrFv7VHbXpwaSsk
G4PuPcO1BOx27tumw7mvn5Ps5We/m5tbahHj5HhWF+OSSmutsy926oM8fHR+7KUXUI2jIKNLUed0
Wwt4oOfzMJP9FqmBgFh45nxHnApiQrOtUWff6mP9QpSb/988sQRQVD+kLvAl1+k1IIl+8ZSf7f2w
DDD/teI1HKXhSZcGbBKXM3u1b7W/PayAT/qaJmjJYCzBF0UIGnzDut9ZJ5BiKPmkjzw1ntCGSZMd
CPHomLaB34yYIrl7J2pPPjbYuoI/Njg2pHuDoNMieFiqFM5VB9ViHq6R849moZ8S8+hyCH27rlOh
WRNgz2winiu15bb73DTe2O50t13Ytlfl/6UpLMlGM0Jc2Qf8/EqeM/jOHDZT37+mlZ09mjUtxRL4
oSph4QpqQCAupirTRKDveQxvdXcM235ak8aYubnGfBBVDO/v0O5jINDczqp1e9MgvSvzXlyDxlMj
yZjcudAuaio0t1IX0dzY0KF5sdqGNjWgpvfT/PMck4BK7TYyA1d39QL+fmzdq+kbwL5DNU3Eyaxy
TRPxlilsCnwE+jhXbShSwngmZfGxBYINR6uiPIWjkeAmZYQ95E7YHIDsQofmqhqwvgrJmdqltcmZ
HtaB1MasPpkefZSRyOA/2HC3QmyU455ximUQInD1Lws9ilnAPFjca7PTpztdgZ5UcAzNN/fGoLt6
dlcaThUCblqSQ52j+QXBXJUgebG+ioNYyGzI0840myZ1O3d1383sAv7j0AprYnFfR6+a/yNqUd3H
NNv5Jlm290K+OXD2AB8003+iriQCghPROQdQceDuvso4CTfVNP40OrlnTlJ3CIlhIy1q+8b68G/r
V/hA8z7cOogMbdrcZnV3N7rtHouFNUuPm9pr5wPCd4OlOXbuZnkN0mHIPD1iRre7aENzuuOF5ofa
4h5kf5t0fG2binylZFSHXh5zDL3BWguDZRs+b76E0Hj0WTfgwYr5cxzHFx7og4YavkQHFnubQxD3
hw3k+F5UQ/3Cz+QYNjuqfun8tLrnJpNxNE4qtMivqPs9i121EupPY6Ot569BRAYslxo4rRtsLjDq
J5HIa+Mh+5QHWNjhQAVqPqRNRnoJNA6rB7dj3+ee6mVeUZRbQpqIUqI8fYh8HfJwbecxe9UE93jB
2aycyldFmff5ZLk5NZlcLeSIMFMyMQ6802T7JLq85/yLMsiD6+CSJ+jtC6x6ICFetr/n0lKi1Q29
nZ5P5EdLyqt2EK2nWWDxTIRmKde8BSuCJhccoybf9rjQy68X0GnnfCZc8AKY/RBLWusXacZri+MJ
dvdrXKz0CmlOxL6DtTiEtw6B2/kqCQDdMwUUcoJnyllXuh5Fz5rJOUpCgIr+6GMlqNmVNEN1ZA09
lzr3KSW/C9fUitLNTwBGqWBm/d7GdBwKG5IXrgh+KjI49lUnfyFNy19mrSlE9JqbBIFLzY1SqwkO
RzJ21gCDSVCifoDP6nY4Lij0lIFGiFQoDM9CgUPJQw1z/d0KHMobJT0SJ4YEhdeULhGBtJUSBySA
vhaNgWdAtaE7xEr8V4KTp7l7mEV1NrAzVzq5JpeXSVCR4SuZ511MYPOQTG1VR84a9UZDyLjwc3n3
Pif6656bQ19ePuKYLhM/sEhpB7qssX49Br3nP6oYAUx2drkv8nn9j2MOzxTJPfAAkpuZ5HWiCKjF
J8p9/hmW6J86KPm+w2UQX83rHYfGgFPNaa0Tp888+Seu3Se+U0ayHBh5RCDnkf7C7X4+NKbU6zWZ
UfceQsyss4FMPi7YzsrK7CQUFDjsksylXC6QHu5cdVSMLa05fRxCe3fxVZTk5BWXGT/o6awIW3JV
HADEK98QyV67GCc9MfHMhrla9qcw141E8GWDkk5YPCKki+NT9AmTOVIquGDrXv3muXVYHmpw9fDb
Pd4gGTF9tilwdvmRl2qo7rzPPgEk3/m2IZkhTGlLZizan8JVV6Penb7iPcvfj/wBhVFs2ndCTExD
d5wGHvuiwwajSgIEjTEOUGk++XYUcoVoaHwOf1pzZtXZYlyTNTQDO6mRQhU1c7VjIEhfD3gkUDWE
M43ddpqSZx2jRbFMfrLJqefaoXG4Ejig8x/oJ65eQ3Y6joPUcouGU3Kktk5j5Rz9/BKcFhMBlnT/
CssAd9AG9NY+Ct9mGXXDGLLqh7k5gtpagoWZldRDzRZUtEKytupzHj1LS9GygcuTIqtWqK7kCmFx
/7pEhTwIGVzyIGnUobtqYuRz/wLc1YPdCCSF1s3pS3zuDNRE00OZGHjX2qyelnXyRcrdb0WS+epJ
Ijm5bO8D5+Liy3ooD7wPhs4qLbCEK/V16i6WvcOCTBdaa0lcq7WZymKY8vnBobJlsmyNGlgFyCys
ynvymItVCT3zhzCjQZWbV22HqlO212jpbkFLO6KMF8n/LXcRRpi3mu8GPxYr9Hbdc5GBBFQGm5oJ
YY4cSwCKJD6YPp9Z1zRZlFQGSLnj+felYEUvDLJ8TtLribdsa/Pa4bdjuVo6a3ctwmh3Rq+oZwVy
2SGVWwaYOs6/GmDX1PIGr8jVKsI6yUfinsZnS4WyyFeNrF3AGvTiquEOwzjSkwbMjGXi/hnR10C+
eYE0Vt7G3zG2jh3OcNnUIGdAF+g5CSv/8OWGN6ysuXYnSOU49eAAFW3biRgycSAzObagw4j7H/ZC
cz5Hbr2NA5l/9h5mHnL3jMJrP3qFqoNBCY+z7hIg8wxIhvZVzvJwETSW/zVXGTaurVqAOeH8mzP0
BuKuXhvStLXXBxYT4WpIHtJR/HKSIUKiW8x7ltFbbdVWPoRIcBPkUWeWvAoJv9uqL8/++E+uN+p1
joHdsU+sXLTfMftbcmYoP+VfsWPrSFbKzujQECIOyKr1uRj9GTJBFVfO6HO6HvRTYTLprnkRM9ru
x+BCniLPvKllhcto1sBWJUEkKaE2Qr7bMXi1PDmv+Mf6SL0koZcp2h9afbbP9q3mXxk+0XQ1hPBZ
tiIK33inizgSuw6vxbe8i7yDk5cuVpEVhf31SyRPPJSaAf4Jh1LBLQhRo4Qj+J6G9y7pM/UYmNoz
8MAY8tHQnFz7jWrPACj1NzsWhipQuj6rW4NZP+IZzYKFkmde0q7Dv6yA7Wq78XveMyvlcsKJUhWy
ug4lqLzD82Jt/kp7Fc2Ca1ZPB+4ghnRKpPpTSiWtbbPqOhdRYZ3yLVHyGPtnzGnOA7H/8JIU/XgP
BC4oMjNPFKxhgfOQRlj+pcvl0+e729oDpybUxcZQX7V2AwagFzu5nmcz70Km8usw9itWi6GhH1Np
e7gCs81OipS1GZr4/SXk8Q6Z7PV/0sjMQN+ZzSkdpvOKY0piIaEYO4C3pQ77X4bk9yWuWJSE1mWI
2+42aRxDPJCdD3wFWQ0XTSb5SiGtxyDqP3yFf4CDlIRSBkrAUWBPIEGPMaRapRpmahK0GBHhZFEe
59jdrBs39Otr875xnPORFdkA/FzxQtx8pGL6s6oRpIeSCUdGb5gVgLVaNZPLAbo6oJoM/VO+M3F3
N5GZWQvSKrvwYsEbUE7goYReNXiVe9fXZNSLGeRJG71orMJ0EZgSasdtqXKrPOyOBaVDb4IXKYZg
FT5PMHWEbBZNv9flJMsl4ywBGQVbN0rZ4/7R/uvm1+mAhIy574vgeNbBOxcd1FzDcqTf+IUA0slg
mKXvN/fgxZhUtp21st++yydSc+DMdBt6GHX7r1CIiH2e4SQXgBhRI00AL8rLp+GMrHwbdWqOXYZF
htRgV5+OTSBpdyXV+Uj8LTomshxFpR4DLxX3HrH5amdux2cJf6px1U0T3Gdjc1EaR439rAk4hY7q
6TqB0i3wd9psuca/8vaRzwFnmHkJXBEGBqDvtYsyCF3p1r2mKOSQ6GfazJwd0cse8Hxs4yosp3qm
ztfjQAkoNXUynzDpaOtw9tLZuz3AMyeqKe8xmHXzeZczjjNWpDICfIgP81Zb50pdm/8hSW4b+78m
uz9ISUQXYx5QP+fuH94DoWIyKNG1qePaXUCeIwhvZ7DhZh0LYl0jgYz61VMc1xiM+YUlc7urSg0C
BE0R9d8v8PlnknJOL9MHbg26UW4Q/EhnV/azSh4KTVhHRgdfqbAzSuNfewjUDYvTIvFj6W5vc+21
FmvxBuYdzXn0MNbqAORc1SQnHUa3fms1MowpkXm2OxyxjUg4/fP9Ez3/x4PWF9HxA53AsxN3MIbP
gNzlFGOpL/Kcx0pDSjCNJ039A30c0Pwk3slK/MWf2te8mzzjJDx0woHr1AkEB5epY1odWk1hUuK8
AlpXmQUQfK3xcYfNibOpWf6HvQwwZTp2xV453MGv/81ukdGx9hivoSshaqKxyDjyY5Q+f7l1BzRF
r5afNOv2dLqG3eM3aXRknG/Auta41g+wRwItyuZ9EvbvA2xLUX8r2mTqmre3til6I8re67VFA6Lp
tx64yTfUzDGpkTEgo61TKVagkbeZ+I11Eq2EI/cy9Crn4rza0jU7trxPkNb6jNrhxQ6mHOtHiJig
eQlUNqq3R7d1r4lLlykBuqkR8vu48ptQaGiEs5pJweLKUXgN93VGXKdLjnf6EXODrr+mG72f8Y6j
qfIcExa/XQkBr6zvVXEKsY/EteVl7gbv9MW7bUOuq57HF7Z9vkOuxYSevsE0VrApYjVUyMdTGxM6
uXRhdrmlEyUYrkuGsffuw3ujhh5FVXyqpjSnGtwXMKqoq11frM1GJ5CpNj6LP/3Z9Sf6yAsCNL42
w3qB61kiQZPeTRsyj4EbC/cA9B+rGTMJuxrC7uFhzqzfuMm52OXscPTr/r0t3zmeVxJbarA0xF8x
7aOYvizONyoAI0eld1FZWBV7ynDinthSDRTfqutw1B5WfOr3EnmqQbMaYECXj6hlb/VPzTucM0xQ
coZOumpJQf+KRaJUNSjxfBaqrSegnW2r+wmMkDiMI1WuLfPLA1sOuM+j0GCc9f59raXm3rJrBpr3
1YXa5R7BIFmfDlf8pL08zeX1e4wIez6wPXiNp1jRCsMwCYklK/EkPXN0T3ic5EDUpYT/AzdektR1
ABz+9RrvQA7cZWr2TLWCqiNfiz3zBKgaPoni/RPd2gbcODheyWW+Y32BVWAU0tT4b5uPrHum4qBg
Acvg9bT/G8vmTR3Hm0+Akp5W4vd2A3G82twvxDXmvEQUTgQGkplq4F2HKgjqU+Iz/JVf0my3xT2K
ytcLDM3vlSNmWodDIi4CJs9UA+o+lsUTM/aHNyq+6Sgw8oEF8pSNPwUVnEZh5VNESs9h0wgfRzcE
oaixsQyqA2qETpdDy4E1RD9vSpLU8CN8U6FJNY++xMRuqqMRRixSb/1V/TwnG0KCNamiZEaSIkdc
+rgWyMqfni1ZneYTiOBQJF1s3YM7OI2kYKNPcwxQD4A4tmz/bZhbGGb9a1Eavl3YAQiObeDiz6vg
ghtwNdKyO9ekontBrTwLtkNhLHfn7UWgNrbkYzPsnmvtTTCMuF8PcHqCfX7Rjsp3JqKMzbIUooTK
LSxWZ9C5yCsfL0CvrqhrwGv+p2Qv/1v48nrZKE7e/JY9e1a8tykcfH50yVCwla+4xrRArSuyzFiG
N8J1aMW9QZd5fZ/YLdnYWvuuU3zmmAfI7XlPWJE9MpQs3+UenJvyLh0Cjkkz1dGTtSdGOmyjYoqc
vIsKlpwrS0MAestLyj/bqqdy/g/2mx55RgNcZOXZqlejndO5S56D+edn9IzP1RNHx+JBtYyxlKrx
uMXGe6JTceKAhCVJT0pdvSchmfzB0QSgxKGcTHOd3JFI/yROde+pVTTHyLknHIaoUdUXPTkA/pLi
3DrypdWpa63FWTVcdhYkhl7wtMUMSleXT7hO5niDQSrd3m2IgjIuZYJOcNNTMaqnL3VPEeVkhEGF
9FmOvBU0tSHRcZHosaZrBwsiU5Xm4KuFDzmMItWf6yQlcumCM4VClHvd7ae95c5lCq+blef8zKjg
AhaCt0UvdAUAOpMaIvPVaGRlmJDpl+M+m5HE2D6P97uPl/43Tp7u+2wh7ypbCRoTMv1WcmythUFL
/hOl4YZRdrzvCmvChRlzzNlojQOnxkptJgpGmj0SGsHxdeL+AZ1yYDDjyKql8l584VuUK1LnlnYX
vAd0EoxS/FzL/UUFHGpvHsOIQZn1DQ0BKFEysBHeXA4nkUgQXQiwDIs1fYWRcn+VX9kQ3plGy8g0
sacLJHsfctMWry0Wv3XBcQtzK+D58lfN09W2IJ2O62FWdmwHt8KW/bWue+GckngR8bIn67cgHJQ1
tmXY7GlCKU6OxKU4aVxuy0OYrcRk+E6CyV4nqGI0q72aHbrfNCWwBvFzx9H7yB/y7rmvU8aENcn6
GvRa0ajhVdUiOWjgljKJDXRx7zyNVMNUOiK5aITDTlJB3rF5AnLpsBZF5KNnCiyAdSM6wXCM/QyW
M/Qqe4EKiNPb0nDExxfafVSCZ/+GtbfTMRBUUkf0uey2FtzJJGqjKffEZw95IuMmY36MxQtU34ey
aRd39ITWJ2DaDtjn0bsfGJW3T0p4X6dyb601ZtrtBn5NKa25LftyXs1KtsPyRksSkwzJEac5VUU4
oyx6MzuUZ/XhaDL9O04Y1MJO1pQfQmV2MlZ/y7E6sycPC6BILF4h4hbsS2Yb0R+94ALEJMPafVAl
rArmJDdk8ukybeGhZZx4UCPQljxsbob3v2C7fAqPDfTiRurAdxcr7KZTiMqoihRDytDnu1YuNvV6
82uZ9G7MA4E5YpW9EhxpAZT0+SbXK4RtuCR2kzX5lYLLKurvFtEXfQXmQCzRQ3AwM6YfYaYbILmz
hzAJKnFqqd1pjQaY5iScyhK0XDESfJ/9pyCLf/VjNAjTQidQ45VDLnbXqu/1QILqw80VgBIZIHDW
Da42dXI0V6Ij1KcMV3+3tM7JTzHFCd/+2FD0LDXt7G3bcCZZUmFj5iPMTWC7cabgLYwcgkHUOMqg
CmYp+lSI8sZAccYnqRddeY/3Ne03ERKhKRIlYs2LEPlVat5uPeL6cugy5k4Wcn3Jf3M6E9H+qTZy
1cYkGzO+BtB+cIpPrq5ZILeBgzBHpiG12JXrS4HtonPRKcPBQxcu/+vxPqw+/7cgApJG03RA1WvU
vFmaazXq4SfewFMFD4t368uKFhnTBOoK+uA6MS5ZZEpVhpzKi+YSFN8FM9bx4DvHpcpq1DcQICwu
oCp9y+60bWLOnOcCOkEOM/+eWrpJzRFr51SwQjbeUYvTyuDLvecEdj8Sk5QvznUc8zpA6MMHUe1d
Tafgvj0bjPC0mZpHvppSSOyTX/qsHMKk1ofCZ1MLo/xjyFQo1hvhCSycHBgvJmGnNVHwG8T6i4n/
xSRf/QV44kxJOTZ7+wzsHSXV5oWbe3rmbyCuqJgfC549JnVTyXshTAgMaBWGPpZfh2teiBVqf9ih
W/Hs4pSU/0rGE+MER7sxuU0IkOZvk+DYB2wqH2k3l7oRy4UkCaZAEXp009npLNWVPzKnJhwsON09
i20JkqREieukzO+m9wXF2HvgXQNoqThQZmsU6yvuJqM8Okk37329Mh5CUs5GWkOslOl8fHpjfslf
MgxYEW05FoQe8S/GZ6tnjH8ktbZtxnWtgDSy6dumhyeEcTl600dpseNMeZpV0EVbd09EzxUrfH0B
XUeOKhRADyo32HYJM4UiyFIqyss5Q0q9g1+k55Ly3587oKJ48FWVmYnGOjFIHdYEdXW+0uCNAU5e
iayq90ePpdAn2FRKSOtHzf/hcuheczZFKdrsqqk3jD/9uOWLHHxjcaNTjX/34aFkE5bwNWNjyqmH
rxBSzN3sEh65g5JyKx36MmpfKgHQ+f4fhzHPgoh6Nkzx2kY2G+wcVPcQ1rVgwCtz4SpGPNwtsDoN
Fj6BSJp2bVUSXNhEDx4iO/vEVSmQG5q+NgeTL5y7i16Fbl8PneBJvTPGUZ/+ft5T5hUss5adt90I
fvH9dTot+LrjqNXyEt0oVsjJLY0YISgiv74AXyLCbvuNqJqw+qkChrLR2lh0xOLDHvqg8tDoCCtc
Q0nuZ5YbHajt92KRG6KX79r87OoDz0s3tq/Tk+gcuCxR40sqV6gYXT9Sa4NcrQAxJ0h0ex2igzLx
9obxm9E3RA9kqTylh1bng9p4+8FqzuW3FINdEJsUo0ziCuzRAPTYGxqNZC2XmXrM76fa48ozt9PR
zCqndm3k4QygWO11yvtzwy3rWMnsi7DBRlcMCqQeHthkszpzoRnHHSBHuyAfJuJFgE/N+Bwj6uPu
+3ePbTjBKp2/Xwqdux1hWIwwThGg6TaazShfZ+xnz5tmO1wv8PZDIdNCVl0yWHgK4DFJ7oJKFoiN
pdRr+gmrbJm4scfWIJOwkR0zHFz9uHgEjieZGYokL44pbdsDhTit0nyYRf6poBKEXyjdePysvfv/
LANUGzbjDURLrHQQz0+cBZKXm7bWct2GWLuul/Ex6u3AR+14EqaNeDjU/bYuemSQREC0V2znF6Sa
u2c1jVHKR9R2qFH0C/7XJM7f+TIbDPfCr4N+We2o7gNrtAZc/B3AEBE4qDKG5dzINU/zIugXKKSi
wvagLh7Xc6SEhhq/vdrZYjEoynHeEBPFX7PfpYahF8wzfzEsJFlbG3fGosrmCu6ra/kIPPms5Z25
TOnoBFaa3iZydC2IPQ0eKcnquC77ZEyRdIGFLNrz//jTnCpvy91Fhib4L1RsHgQtQMlUo+2RqXBa
Lo3/3Lq1T2iqS3P98oP6KsYxk7aJG5el9cUGGnflClmleigm4CW0ZRkpv+x7qqyXfkeWlupPSlC+
K2F3b/pzluo2eutJlL3Wi+dntZOtHqvj9SCM4oC4E7Ms+CliPqnENDX83jhh7ixxAGbZor9aKLIp
AOb/hAH37MW16enVzyQ70lWGf7+nEDeP5d5g0olZSSQp45OBqbTmKd9t6UiqvBlcEwlxASJOgr5N
Wwj23LwmTAp6WVjZ6ZHvh03fnHwlP9+ZKyMwz6gcmd4laBLSKOhaHpHAKYNMAR2ZDSE1nwYFQXr1
mJ+/uuqWzqn5R+qjiDF+dIkDg4f6zs3eL/2TBoJxyQ/djtTiwochDWAvnr19dCVSevd+REUb9z8P
Y05fzQvr3N1fqI51WT69GyTU1xKy09aWKjKvvFn0Do6Do/ILTe0jqhwPotaNKbY4MweUpUWpXC2s
B/6o/+oDFOUHsFTwVpThwl4/pBh0upHBETQ1jd6qrrz7O69RW9n8D/wVqyPatYH6wUbHCGNTeysY
or0QwScQFpvQK73AYWZCZhTx76AdjDZHcVrove8LEKcMFt/DfW6IaSWlqzmKW9ibtUBYWIn3bKim
ZMuXoe8ve2+2wWV7dpA2uuca8FNl9H4pTvt6L7pxwHIsbfpR7p5K5SeefsRIGVj6K1kcTFFJD6Py
p/TnxKTNjNW9IY5v2n5zc2raqbrqrzsatEVItgrDPdvfzBrMJQPJGD20jBg2Q1hKj4m5NKmt970b
c++NCiidNN+AqfAHO1wleO1EWeavosuXNcmH8Lte46LrK/IB43grEHkwtjht/4bCUA1k3ls+O5Bv
catTVnFUVktVu/aFjVHLD4Igret11m+HX6PHGVax3gETxmjUkWfI2NxO8eDRqFBKPvxrrnre2Hh6
otTSVnKRmqlxXBFEf/cSp1FXPfoYI0z3A0XrWVS9ZQ38fYGgJdW++ZYEEvKNJZPkrm2tWuMqYuob
LeX/U/8w+A3sonWdAvBky7qnZm6IUsqFn+O0F+zkP/Y1AzjsLlvhOXnbNV/TcWAA0EXgDcaBDfMM
KrGnPvu0isn+CjlWMDHpzopSzf+sZ93tDnQMdmVm5IXusyc+dceui+B3DyrZEnlKcDhoPIeW1rUT
Oe9E7yPiOx93ifxWGCnVHndtzmlWfW8Jk5hs35lJUuySuRz61S+HZfk3BEvVQn5Cyk2I0+ugsHlw
fArq76YRtWpHV+hKjgSZyp6q/uYv7M0GOJT00cYJ5NPVkUX2vNQREIQxsG5LowIgRuLggp1gj6Zu
qMznaC6Q4q3if8ATtke0FMNC5/NT0Js0jHwUgiQ9Rrpc2UJIIbgJCyndrHse0al3jhOXm/FwRCUU
3Sv+v+jcrD77duuAx1G38pdyt1Ge6y7GOyC67I2xUOVkx0I1/ybjOiEw9PFteJxhCpf8mAikj7sd
/PyKJIY91bvDfLHpcwXa7ZuIL5dSWzoHIoJ/KBRklpY1i/Fj//ZGldcArHPFqkxj7BEmadOmxSN7
XCa8ZSGkNhjQ3qzrxj5M6wcnoGHxlp81U5JwIj6pjOZrc+Ia1mz/AKD9GZWS9n1foArOcqzWL4SS
TiPrNJHtl9uE0yUPzRpY2B22K9ZdBceLOOXfHIrpwhlJZgBbxfrdN6YXe1r47YeQz4dT7axEtyXX
+d3qvhhlo8+RMq15y54LwP/yguhOMXNhloUK1zy3lcA5P9+tD6UCjtuO//FiC1W0xMl0NLvYHwXM
U3hiFtp4dDmTIKE+lccgoIEiePXpzMiF6jyrIF6H++5+Ntg/j+Agw85Kr6ufCijLeNdV65p6Y5tk
AbHc/PZfXX2l1tYXE942XXqgjBuC9A2Iq3WQqDE+uD8Py/rE9TJzRNAOAijgcMebxTEsPFkgvWbr
o5EBJey+XW0+apAWeCSuVLIQQ9MMDr2zSzNVjjtskNzmrw6Y2BUpGMJuFHz6GFCmYsM5XGV+L+zD
9WwiqwKQWDakryb3cfl1gyF3lxuEdKQJZC6Mj5/TRDBrYuLOxBcTN84wW6gocqVXGkk2ImWJu7sx
kOaNukmeGEpfc6LPHnrcLteTa/pFqkwBybVtm2GNxA2uhenbWFYsHf6WUYAX0GjgUuEhECv0U39m
4vmtuD9t37oXj7Pr5k3cFQ8Ovqu37jsLCXHDbCjOQE+EQ6BWWeGgPEVq0vZ/qoaW66mHY0YFnssM
zicPR4WsS5vgg4zGK0Y6bRmNpEZPcUQC4N5BFZsfNXse+ur4fJ5VbJ1bvrhr8AvDNBzqbTPnwaAx
OdbtRyR1sOUAgcUr7tjqPcta99UcoPIKhLQi348Tollf7o5jNY/q5Y3Pv2H8IauhatEntkYYyNB+
qXAkIj3UUJXt5IzJYQZq7kog2AwB3Iuu9HplolyVXRb06A87sRvJTTXpL9aliL4C7ib3tCT/F+qQ
PjkNJ5W4XpYBwxjEZUHyLlWLROjW0VMj66v2dQ/P05HH83hBaOcJU/r+udOqq8g8lM+NzNNMKgIg
hBybg1gKHzsn8oAxs7e//qaLrrvYuf+343Rgainq4IERm8SoA0eY/ly/YCFjby0R9QbWA8pBAsBl
YPU8TSCWOCTeJ1afLL3miFHJzmsU+uPfyYh4pZD9hns9ajni27j7TY+hXZN3/+JHjVCgZjZYK95n
JiFGDsBgOsssKGP3TuGaArvGx+ZSrfzeov81iLe+BkgnuMi8yfG2i/YHHeAsSyCZ72GpvSC/I3ua
NSyXsjZQXkDkIWWc9nuXHHBevprOKxgFgtlDjaeXBLGN1ulPynhL+WS4YSUAWbT8fQ2As1yLJtH2
UC4Fqqn0ZN+zN8d9XSyE1Z5T9CgIaNovSySwyxRtsLztaakmYJS+SWsA0AYtIfXKxMR1LPY5e/UJ
HaX5bdB5P2QswF2tmDDAF/GCi9CBfhA9Kokomg2qXzXZyL8KCEv2yktgkJU4PyTGi8bOVo5fDH01
WpBFi96uqUs+3rh+vFyXa8aBuCBtf0GvxZ0TubH3LUBlb7n+taXMSuScvRFrTNIXqBhMJJP4uiTV
PaAerpc0gPy3EMzu6MsZ6Z1TrTEV7CqVh2++GsIDm0fgj1yFjA02dZw1p3RchOmgE+b1KGCnS8c2
M7xlZG6QZWtSnMqAYV96tgjE+XCHYlrwXOTJ9hzF85smk9I8MqMRpLbkFTZxqutztv573Y1oIs7u
B12yhaRMUN0SicFl77jp0Fy08EI5xQE8kLAethrcvxgn7048wwNUwUbQL1rHuSpAQWjfixYkLOrX
vDi98CGX+6ujuu7kbsRWF2uPX/XpnL53sViIBNli0nGiFpn6WOGSTdrOiLv7MSdLd3cv7wEPWCsL
ufF9Li843Zu0bZxHgKPTi6pDzOlE99c+wadYCYIH2x5387XKdNJ6Sz/XR1KLzLadP4QHL7THn/F3
tbBx7k8yeHZ+KNmoew34IOJ7BZHzjJUBk2ezqFcRHFm3W9AhfpgMbI1qcGhs+oyQ54+ZwV8zkA7F
+ANvIaPmF4cg+nJrP7VtCfD+9TEFR/wSfRIqqRBZX8pXro1dVfbKZ6Rs9VYFEm5tzO3CxxwDobAh
adoc0S/c6tssSIxvOGb4m3mzMBUZM1DvjbdaBXS9EhrxN5C0x9tvlJzTkQKY+TfZKcbsL30flznn
rpMPMxycFyMqQXGmk2KpbORlBhSHj5T8ihNEdEP9wzQoqhp18DXuH6Fhbu75LFE94Hguw+wF4aId
RMwEITpSbgswbiRmgSxz2MXyP611wOZD41QkMOtx/muSBcBDFzuZZiZynpbNU6jLHarrUdLQI0VG
7GBZs6R9hXFqFbfqh8Tctss7tYuJYS5UTA217nMRULqzly556AzEgrwuy91XSbYFa3j8eOaFOLbK
fnMGxrLdPumQE+E56Bu9qqUT/e6pKLKHxqk3uzv8Ncj8euc2O4TGNvmr+QwUCQDXPUni5PMFjmQp
yQTWaVQVZ/XkPewlAfoOgaiA/U1uDffmPdbCgGM3HKnc9t3JWwDEdQWwif0K/auDDrP9slQfURr+
CcYdSfsfeyu/ubeIUOtPglTuyZ7xWEWEeKbAvJh9XZ5C/4A77TAngxhG4z8Nhf9lNlor4vp6Dzl4
xSEWJf4E0F3KB9fndbxRCPvVPaMM1NtyrNSDqadj/TB3RJ3FlXaX/saMNxRa/4plqFmInB6V0cY9
v0gtSZYXE4IjWBz2zD8iCScyMP1iTTv/iXU6cENZJ6ApUs9vcQ4TYdLjvVg6vBr6tpvZChdOTYIZ
tEYaTixu8Tv22kNlnqkOwYtbrRr1ZsLLH+oVhY6iP3Ftp9zstJ9SRYUIC2k81SZZVleZpusM1WEe
tUSKq5TS6PLp35HKvIs9NNWXVHd1wIAn1qRFxvOFPsykrMGlMdgtRkG25LM17vnkh/Z4mSCaHkdd
iRPir0CXdxKqRXsz+fcPQbJe9d2iv3rqN47nAYjE2bdXLAIh2mOmgqOceu6ISXIpE2f4WmebD3b3
cme1hzULZfgxo+JBWBXxdtHcSbTZw6VmuL3LjvDPBw7u/9/rGYIMvRbWlefw8H5WvMbeBI4hpXS9
9vlmfluWRuVE2NnFBMyTwqwRUVgHqDvwfNR3lqrNAXM8/7I6SB05ovnwbpWinUq0ucpGZVqcRsTe
LtNkv5+DgGypEAzDIkjm9frCGMeALbsA9+p/aEvPtDZnqkIzK0bsecJWhmpNC7LFSgzPzMhgghBO
LxvTndPU2svhHKuybGzE6tb9t9277hGKn9J8JGNs1FCTGt5HbdXd1cc3X6hN4iamYLqB6gDDL+uR
fk7tSlndwENuc91jUYTDanei11ZX7LJfOh9g/AX2fIpxzmO6ym5Pt6X4EKLBAkKKHEkzXq4WuWEt
nYNSPIKELJ0kAeZtd1a3pyBQh94LR6D7T7MenpVxK20BTSiXbXTzMteK1bZZm0iZuCdSTv41XFV1
8fG9Ho89yL+Npg5lNweVw5ICz+uSMvbXEUuA35QkFEfC0Py39Nnpd12Lhi6aIxEwEn0yYTEdh6xs
TLfaOFvInZ8eWG2xYsbRRu2OU7nYzLEaVVYjY4Mt8jd1nb7sFuCrCtU9kPhKeCvYryQ+S4EFhOmF
fp1ENOYKdvrPwem3Pzsa1yn1ZhWADDuNOy7vrW4yYJzNrJb2w3L+AsKKYqbC8JQgi6WmffcE/8mF
dZlXt+orgRZzVXusFRul5ukAD3ACGRuGG9EkkzYpjJs8Uo7V+NVzVXO8xckwRV4hGtyYm7BFCIJP
11IyUmShNP5PsBNVVURWKqOq2Q1y4WJpEpMfChjXLWMQGcQetWqmgNzc3oYwIhzeEpMuU1py4wqu
F59Ub+4GIn7U6JSFsPJyO5+GMGGeR9ELvLL5rfk3hf3l+enVBu0plnCEw8XdxoZxUAkg479i7g5z
iGSyeEv4ZZqjVXR/lI7kWZU8ns/4lxepDwXYwrHrGnbsnPc284v5tPCa7QDy9ouzdoLVuU+SG2z2
G2GbnZNU6XOI+UyYqHeDV+IZpQb56fW5A2z4bd63kAiBHTQOL50yZTnrBp/lUtYt68zxdUgqO7US
vCKo1iDPaluez2K13mAbygb+PyliKv6ZfNQkLqqzwHgMzwIC4ifi7dEOC0fJn7xPRtKycJRPzYmi
5r4l8S5ZFRAjJFh5Ycgvg+ZUEmC4QdL2P5sXiZP3iPWaXdkQ5zw7Gwjqy1djV4nWqXVRBLdOCw+m
qSVyg2wVCyZHWmEobzMp0a5Z6reLNQVNEMXtXmAnQKuCrdlnE9pDfl2b4Ykjta/GdNROPEw9Pgb8
i4guAVbzRuFTg64R16QaSuEj39vvhuQnPsvx8sHGv/Jt3s2OKrmRp6uH/5G+Hk9qBXH/xs7FHkPG
tTU++sBsYw7jQNenhhKRqffTVVc3WlnvSjznNS4oFycfYZAclAxhPTwhmsPH7bIJtypkU8sVK5Yk
RAo50MY9KqZkMDUIxmMSb8kZmrzLhop66iEQ+2FzD68tV5HdLsDkcCMona+vHzztvAOnSIMzcq3k
ZdqvQvHyVzqHtYU/Z5M/HBy4t+yw+vltqKEqSftmZZ27MidaYLWY5X73HkN0yEqmKhgc8jNp1FOj
aoi7SjEvFzh4GsiLK4z9dIX6ePHm3n2tQhU2ABPgZpfDpj7Jt0KTvftCRd2YfMF7BsaGdXKrBQkp
ZpYysZ6wk86Dwq1oo1+pYQyDPN24GD+Y9GoO+m65G2rJxbcpah8f3vkFp2jmlsYUB5VfolobDwQi
umlRMjruM1q+nWe4Vr1BLSwHpt63RxzVrTMhAJd2WiWovpJDZW48nz0MLF56Tv8i+O3BRVU3mNCH
CUq9f4l3q/qN1i4N8/DwZurbiEmiGIeEJPmz+2bN4KjUYevKylf7tHBTRGtVSDm5pj3Y8xdUva5r
DPZFTJishPRYbF3/xoiMBr28Ppaaf969EXkE4gCevbgDQFF74C4uyVZz4ZX74fMSExn0g2pQeZPX
5vmqTfVYhIqofGE8m+1AjTjvAZLaffZ8yjVCdXEq5pKSv3sN1tjCd6KulVY1ZZZ/bVFZhe5U++y2
3ekhLzf5SKxX9xUR8Q9jN75XQc7hE3KcBDZX7TTkiZtHY5oyzlfppziT1nrMyr+deS17AyKOUYP+
UQXCo0k8ouoKFpuGdURYFdJNJgs0mVazEoZE9laDNxFW4AxqeYQhag5PvIrFht2eDdfXQWgX+ya3
g7NMz1MWaDE2P6FJ21oLilldxER0AjBNnzTXik0q3l+nMe7qWkBnUutMY1joto8tfMJq/S8HGl+t
U45YApniaSxpLq51kWkMVZ7aOjixURzHU5mC4Wi05CY4aWFPJci4wkjNDGrSu99JmrEpbvMV4crp
OE2+9ZpJ3N7VHRZxHGvE+yEi8wYpJoczeLb2wTQAbKRel56OQQc85VELQ+lzuYuAdCkdzCbDhoCX
gccLgvGuWe5lbTxLOexX0ZTLmFnFT9tBXIrJ8Lh+xGR7h/UCKZAiWBbnk1zQtXoRio3d7VdIDhYS
NDpOCXz1qM+dnV5dJNdvMEBUnxYO9Pyd2UHemtNRk+zaWqsT/mz9I9eBaPd4LZZpJPjOXILrwp1H
B37hGOnrGlBafNmn0s0Tw3T86u1Vk8wEQA2DEiclMgNdR2OpYX2ZFuufHdEMGbidaDqLz3/wyZns
9ZMZtnocivTCcSluObwb8QLpIjBnztUCrGUYplwO+BW8o8iUP5n8LBwydimdtn1P0ZrzE7FzN/DJ
ZyUx+8sXpWmBS5YFVsE/xKxJRSBi1EJLn3Vj/gSVIkJ8c0V8eC9H9Li7WMDCrUDxcJPpb18sinoB
e0PzcBdwrGfOBXQ/EfzZvibMDMewYRkkdthPDqDcRZkzqnEgy7izpDZlzQaAFJFIM6FquTBq6knA
PEqHx1xjHm4BqroYzQ1nJrAPp4LyiRs0Kvg7wDBfosNG9zO2PQ29AtY0inCDqar93mJTWzqhP1yy
q4Uf52fR2igb4HJXu1D5lCVK6e/kEwsfRyYupapc5bzQwUAkO2277AE70AINDvmJq+6sYZTB36ef
RdX23bWULnwOwTWEm4/yJLcEiSXHcSRreGf/xVIi6v7AMUgTzJJ+S0vJaVaxCk+1NhQ+cVxHeKYZ
YiOr03KDlpBScFFxr6XQ0qO8FZTpaL+oYRwyCO0k/M2QbKAOEiYvtlHsR4CtJdmXxkHTXYrx3q4Y
s9EwNj8Quwou0mrtjtFjYcNAjBp+jaWMG6ti/Wl3jr0PAcqvAxjc/Z0+4TBwNCrsJ05HhCB6Xx71
Ff+z1KThPrE2fS7uFN080yKC1qZI5qoyOyJCzF6pDfMPMAWMRznJMKjz+m2x8+/qruogLyFMrGdq
Ik7Dn/NNlgSqUdr2tlfSk8va6r6eugz2WyBUpkHvByuJuovz+iQH+MYCb2t4JY7I4wzOldPSQcdy
m/1fS6ixuyCDOjogKIO7MYwKoGA0E9AHLPH+sbIZz2L0SQeLifrrLpbb1OQ34fh03XRB43vArb7r
u0bXqtuRVjcGD9YGqXFYPnqW5Xeq4aaVzMhpJ3utP9VolsL2VDwU34NdE99QSP3SJZROtXGJkp0x
BTPPEK+X0KZVnrALHdSw6sltNOq5xbPsVoAdHt4Q5d2WMK0+JIChMn8XvuWwEoCT11MkiZYhofC6
j2v5ikLYHhEOSBXrtjxDhJ71MCzIgScNOe22OEu7oUpSyHjAij7ijIBf9bCE0AB1FwCKSDJ+KIyo
9MV/S//+3kMF1L208aThKslPP8nStDT+1JYA87PSh+IhFgZa7C047+R5PPIYdcwadIXYAWNGSYgG
+jVUFbIyk2ZXxPl6IEzIbkdeBeG0MJIsSrjX1faugBLzK+wu0T0k2f+D0FebM2v6oKmXos9mWDyI
7D9ydEEQ0Vm63nH95+jkXY5JNMOtdWvEo03LRfSmz6lRa8sjYXI0FkMod1L6fnF6c2x1KEG/r5JR
8ETNEFATxQVuzgdh7x+RLaf1m0mLQ10/UdjxKy2qHxbNaDHKY58yybfktC3CpijmPdX6PRat3hwI
qMxiwxpxoSgbLvUV3w3Lf5yNTmcii7IDeEROE7xXA/kWYMVG8S1kdHsao7GvGcy236wsw6CfNLuH
Qh6y2Th+vQvQdZO9Hv4RSMKxvGxu9ZSlj9v2hdCJDUPglORUS5Unz5zxTMErH40LEnF4poZOfnwd
5N/x1RQOW7GI49YX6chiGQI94aoVY7zrfJLHenAIOe0Mh5k0OLJKeyxqZRWqbgwYp5CepWuaMlpj
w07XEKSqVmg47jduCxpPklhxpdEWaIKP7wWRA9tuxpTr4wT2Dhfj1/rXY6GOfHLD6zH4+mbZ+nYN
Zf3kiRB0t6WyKao+VtmMAWea1T8zuT/iwdOWDuwbQfZzwSAnlYJERsppoX/xLfpP5/HGI4TvFa2c
ZxSrdWIoRKNSuZ+UixxPIVESq+F1kZwIl2s6jPjK/CUw4AYZSgxq7ImdpMerikzBmNS40z0/lVYF
SG3fXayJWfDoYvpkQCwNX7WXzNksTBU+I810lbw0H/KSD+OH4yqnviIpzn3JZtE7ESDYz3XJcoKN
mWf9JxXnmsuDOasPsrtK6jnR+Wyrvt1hw9eYUc0CDyK7rxsTYjcwZubrDNDx48GeHmKdHN3j2Tdz
oxoRCobWgIOmvv2oU9oRGQroNvQ56Ben5ZqVqkUw3PCBjVMEzOv5lw6Hz7S5W+Jz58QCTeZSwAmu
u2DE5dA6iFP+tGEalzjUnWH1XVPcPP+V7/q7pJTPOiGoQW1CgLWdB19b3AtRTULTf7brdLrETlsq
51Gio1Q3203K02/EYda20fQuSjugYrOb1wThJkiRVE4/E76ByF3Xjrnr5HJ8TU00FTsTyNTJLebp
VZibkrskko7K4MNvFiGJkwv4tECrBsNpP5DkapZMsjvN8uqLX7rSFrk8+nBEA9N++eb/0tnXjoJT
OIapZG9W7ILkiLPEv6uhU+CQU0wtgT5vMEKGwJK8sqIxoYgLI0lBsyjCzWFtjlJqYaq+wGJAo/yi
M89UvKytBFZ8yWBQkMqzkGYPWDEVZV5BisBquZDyFBf+XV25Rk0EL2rff6feGMumQcmjoNO2GGv1
VGJSVGxyRlNmBrGwV4mkIJLCNaUzCiKdocFLnCahvKxdNPz0yGZIqgZZqxwaFtu5KyGn1uscmpDd
9JJ/lgTEueT7hjs++iX0+kp7grJkHw931R+Nao25DGgV9Tq0X42wdP+aN0YETJ5ugY87UZYmJLj1
UiBrPBjwvnM347MFz4T5qaeT/yAEyALqsf3p/qvn9AFL/AiHTAzviiMg53Cv9/+lGA7dYsPRQeWq
t25AcANG4J9Yi2A6xxh0vwGXM845/g6uBombAmUjzfZlDgaTcpf4UQ3VRiZcT/UlON/c1s0MwdkX
fiZ3hHES6FEuRzS/14aaBcjoVpjM7o6219vZXigAkcXZGNsWVa+WLjLyjFb3TR2myf6RXHRmtIqp
oBp2ZwmLktZe4a8UzqwA/uxREF34FzWZmlLVqA0ajrwZrA59DUv9Gh/IpQtG/VKCsrSV1vY0vjUI
zJymeXsl7OUJGt0zflQizQ+JlD+ywkgGH6sNH7pR/2N65TIZtEy6xs90M/RYcztxKgdTskjK2MZQ
NlZ3Wp7/kLL2dK7c8qUjiuua90hxdR6LIyxOoF++CgwH8eKBJYVC0dVY3JV4lrHK+X4bxA0KWZou
ona1cdyhud0ltZ552FyM7H6Y5SOoUxXUE7OEfL8sI44b/9sH8Qb+BukNf0qccMoZ7zHKxRnA8s4w
tE3puKcZTlcScVYw2phxcZhRWfs2VEZAYuu9NUWulOM4bhU5pG8LeuWZ4+giSwQtl3yonPLh3614
WOs8vjR7DG9TwMGSwlMqEDZnPeAetYACd/D26r7raKBqaakrT2alJHYmoWhun9GHebE3R4PnU9c/
ScxThVtG3IA8qmTqnTZGEFWRt4Uew+9Hr9TzFVzqY/bVUxd1fH1Xs7GBVP0IrXln+XSMdHgGPpzq
/e3AgKWBztTI0fRqASlGeqZcoSR+ZA27ZOvEMrIob3jAhSoC+QGNqPzNpeZoAyP/As7BEGvGFnNi
GbmRbya/4q+c/rmknWAL4VViz9xmAuq1IL98wLaxy6lIfIFXvCPjtpRZqmye4RAShpHhhsaRx5d2
AKWMCId3OBvPoCt07YszEwgiUzzaxwaw76/+dcs9gX1Y7SzW+lN1+42GfGh0lx6VT/KsVlAM729d
uv6AASs9q+D4ANb3Ug4hYtBdfwJdD86iFRAW8gTUW3bniKemAvlY7YMQQAiItKuFG/wuk8v0vFV0
gPd5pm7ESAuWoWkFly6ozoN9kuQg7rKXs0FXAB9jXfMXjK4648/eOe3/G24P7x8PqmT1NhHohT1j
we2E0gstMzfuprvEbpvQQ/F4ZFmcfGNLcpHcJ2oKpRShFsnjXZY3lRuGCsBBjvz1eAaBrlsYJ/HH
UgqHCkUGfio7tEsRqS8Ge3DRxIFjHg66+2SEQ33T2Sf98QIG6hjJWxicqjnjW9r0YY863tEkGIlI
Q1tlVfCMKT9AEjZklyFa6SaqFTNvYcBTfL2umXZAZSr0SYTE4hivt6q7iqln7Zw6zbjNoLmA8+D6
AA8SIF5Rvz5nq2QJX2zY0DBlcEu/TOFPsnbrml0sGYWomXtr2Gpei3WTKBQpLKdSXi2XZZcnAhn1
0O/0pZtehHaLEY84O9GRY7VBrYnqfXmov7XxSDGYEFwdumndkJUs4FA66f3duMU4zy28wCkp7rsa
Xh1+wER6iF8/AtNzjGr2MylLqTqOxMpsWiIBKexXDtFH8s54hDOVar1+DqQ5anFCO2IWqUJUDxmg
x7UJNZOpxs8W10WOitrhzNIfLbs2DL7nksZyBQZlzpWALr6gyQC5dOiwqqkQxeEXl7J3PIfKpe5g
645rygaB/c+biP7pKfFYsFdTiLKfvpM6r7/qaZWiKjCWX51JFMX5Ud/kkOmyK1U8NNg4RI//0559
4jGauHoWEP2Rj1LISFDZTs9TthD2ApW801QJcDKV1lgSLNLeok8NC1wvxDDw2UQGIxj1M4SkznJR
5bBvCdoOsW4d7NmSGDAsk3YAqFwkj5V1P04BZ4fnKbTTIQaoRDdBghq5T62QlMaGIByq/z+fTYq/
W51efSFhze4ab5GqC83zSCwIOdb2BIUCm7crJK7B58ohsotsSqSa5JvNgIKivh8MBKy8PqyDhCcr
kc9OK+GFFHqiEtD3MNgSEyXMaDBZmiI9hIIAj2wfcjRfoeeMOyNEGQA0vawedcrXRzitaz1IwDKc
vVek7Wwyu/rTeAxSDit2sMNC6T1MTcxHrsMkiC/HmO/R1QbYMsvz//zgTjm0sq/3QlaZ0Hnp13WV
U6f8G/3lfFcIxJ8UbD+X24L/U4cvI+neQf3OJ7oRIAgIeqsh3zW1ym0QvORE77vBhjwvHPX0vjcu
kY1JzXRxqKsCxqRRpjcsN16/fwMWP5a+BVPqqe0/o87k5GhIUPGswAD7OuCW6GB/p6F6NbRJlnTj
wfsNa5vqR1LOnjjBA6YTyWnqrY9J7zyN9Uu9w+dep22nSoHPmwpI0phyckorsrc1v0+Ycuo6XU8K
fGyZqwqjFGsBeuYKmG0nOyEw1PKSy6yEB4IQXIpIeYQctRlyfQxjQX/afwCyaJZATQOdvAWnVG63
btvOvByz2xQm62YuRjA7xpBqTV3PEn9z4wiN7IgvUNiOCb8KACoFcBK6XWZfEC/Mgor3mNt/DGAM
/oBDslpEdnmOS8OoWL5w2wgnKB9TkOYv6vPUCMNvkXb8jvL4HTh0p7rWa/NGzlnas/lLGN+cRFfY
P/F7aYbljnG+0xOKBzzngRvxhhi9ydOUJGYsyVqQbTiYqGy20S6Bvp5J8BbLVEYTv/wRnVHAeg//
2G4L3v5pw5enGTkyh3/Rah54EFU4iyOfVg9gIftW8GJNJnA1hpqEPmgOWQehm+8oae1rwK2ws2v1
gEQRmLdbW4A8wdn72S1P0JvHYCP202VzGfWUhAQLJ3R4eyRXamLy/utPPy4UAsFwvNn5dkiiP/Tr
RcbV0yjb7JJvQ2ICR5Ce6BCJ5DKQisHvK/0Pby/u+OGTzoXSXahde8IrV0gAYcFYOV+UZqYgCkC7
ZMqMRyDwq6k44Rj7tDKMERSTr6cHLOT2pQrZQeyRr0mg0uDqBXj9WL6wZqQYZe8tqCeRqMnAbvbe
sUmheYCVmNo82+2lokYHiolwl1ELeWvxXX7oBi/M6DE/TMPtxzSG8RJ6SaL14DZ1tqVhxNtU44RC
kuvZQA0lh3Go2pFL8XGqbyV+kDxISuRsKT2PMJ2KLiRK0KSTdqTuw77jeab8T9B9RKaO5JpWvlnG
THRq28nX6xnxnp+4QOx7aY1AZK0HXQu8W3iojFqe0AewA39DbNByoVibRaBJfKJJbTW57o5kCGqo
nNIqwpK3hSIOYs10OwTKV4Msa0lgd4ibE6XwqCPixpF35OViMC1Z8iLxseatjJjyRS2nadvNm34v
JeK0tq/5OE/1RXa7KpvhprZ6KM4U42uy91V2TWIhXzXbuxEEailGVU/hPvZ6KJ1YSp9Dv3rPKIjG
/yvaS6C/3YewMrmrkJwmbN3krlsqhH65qJ6JdelSjl3l3vK6/Rn7jxyrwhZ1lZfDb8JknnjnIKb9
sB1PekdG9zX/xfOTyZAVDT/7eCzi+SoKZGF8wf+EXXMetLSyDNXoBfdOXq3umwam0WBtHWZUsO9w
bZ8pC8l4jkYRmNzKGN1E8cOpBJCYeSG3NbsIh5zZjjwCi9mYORDwYKcKNUFglA6ja7pGemeco949
bUcj03xHabpJ16qvAWC/s+zsnjx5tYkmip95/vbaSy8gND8axliaQ3Zu0fV+D2r05s0SMtHeqsj8
3rsR3LD8DoAs1xu5qbahNn8Ik5umW2qPmAJcEkKO2F9BJXSwgWbUIi886s5WcZtA54cfarez79Ro
nvWN4s6IKGDAMxcqkxuwbcoPhfMefwFpxretGAkgWbxzQ72AT11asrscyJTV43bh73IdthNSP1+L
0H40ZCWh/IZjQYWfcXtHG4dShBlnNCquvnAgRyo6nX9AnrIePJrYe0PmSssWyaOamt7YD9UcJe6e
FDxM+sBMDVYB+kpPAj6NR3iQz+wve/8oA0irwTy22TlyvdN60nV2o94Tjy7v7R33n9IUe2ITsM6I
0sMLfUpaXLHv5W/9s2g1EDWk32F57O1X6uLlREYYyyRRPirf6hVRS8LjZhwVWUgXUt+R72Qt2ZKf
BmLiX3Pqmc2/zfo6FT7JZHIxts8j06GlkHnzxusSpN0JS2SYYb5IDJu45f8Ylm6uJ52v1+5bZlmR
ANcXSn0FZhWy5r9DaEUIGZ1nUOPJV7kqLRG94Y0H3V9ZK0ePciKSK7J3n/EhGwAmw+gpS4ENwPio
cO6a6SXT/RR+KOg40QIcWk9zdZdpyl7wAgKGEORXfZdTTDzLoLm8orbtCUmEm+ghe9Brs4W1mANe
gObEnPoacX0Hk1i0LR3ME8k4GdUveWKoCHRfl2Xvf1zJlALrwGCevxdwV1E9U6QTQxR7r8/YiJEd
/W5wyIEO1qHsp+0/ShR1Ku0aAYGV0YuBV3mPAACGMOYf7N2TNvRgb2vtjg+FEX9Gq1JvkTfeMVDa
tQNHi/C4a214X1cgWtzlK71BUo5YKt5kREle4Xl3BV2vVvHsoevhU/WUAIOt0lbM0wNMAYTfdzCm
19H7KigVcsmNPbLvdce4t+1VR3tjXSuy64Z60G3gzLSZUJpsnSA1WoGugQr8aIeV8wqfjkt0h0f9
pJU0KUwK5S+v1Q+0+SzETUj7dmi27SLVmaRGAGW+WANXlH68Gy9tFVLCMgRNCNp5ipU94AXXOKMa
2DhSOo5SaNCyMXTpYsqSMbNBv9X7tWaeKYYmWOwGE9wUPQwtkl+CkpEcOzXQTACMovdl4j9dvfxH
vwbjAyp0IPT3X7JGZkAvWCEycAfqfaXugjz3YsnnEzJWcb4ZNw12R1ZYi353OuyR4cjgsgzpKemP
Hpt6TCk0xgt+uSdKNiydKd08aZy9FxI9/kACqahW//ltYLFwkLi6BYgkSzQ0rL73NDmDpD48dXAp
SA1sOGII/1BD+oV7Dd+giwzvqHAW3hu5PpjNLtTQMUaFFzwg03xpsVRJJgW8UbECFlFq/Qkxmmw6
LxBzD3lhmVWeKuLyryyDPhapa9TJJzj9qsxcgPvrn90H+pGTrzfo8LyRrEedImMdpMLe924OVCLE
MQwD3dlg/ssSnEwBTPean6gSCUX6WMSm5F+7o0pJt57QikbWtgeuOqqLZMneRcnqLoMfhXBaHC/7
js2eIo86qMC4msAaLTkffU/z+3wKBvzesd6XI6WdaMTGwXHRkrI1vnK6RNWtBq+wme1PTh4omh7z
BsNzKrt/ktNXOR2VQMkhkNHhuC1SVlTWWfiHIBzkOBpZXhOVvdCHLpPAUMdkyyLwNexdW2cjfSvf
Z2ep9FCxG0NqkdpYEAy0U9ASZklwkTAzAtKc/d4EP548VBGylsJU1My+BNkLXN29HrDtTNh1e0az
0JLpJFROz65Z3eER6KapKiTDYOB//fw5DuYtp+tIl95nZgX7TFRfh8jV4Uow2O+EnVxZfrODe1Ex
NTa8XOOMto2AzH8TS1+u0DY3wj38NyjvKJwCOC/Narn89q8EJzcM6CqonQZ9otJcAhEWr9XPF3LW
Bidwuhhoq/87OunUq7MTyQP5+kh3UaCzot0FU6aphOY6nCCx9bAyQVsBUIBKl5hAz/3+b7tpdqTW
uZxQpDcGJNT0wgfbxVG+x+MB33/7gZ0uFKQIcxKJZyhPBAkJ506q/mTPyjSWsSrJiT0IYSv8x+nX
vjpsmYv6LTIdg6GMwIUcS20y64HFqh70cPy1FAxcTSyt/w3mQTpw5RxxxZPb2pcJdBi5ZL+2Ru0U
QM5z9vr7d+MS8AYn1Wh+KdQwyfF6NRNyd/XZraezkt1KKq4/1+0v2QWHfxv/KOYeuQIxkJN5Qxcu
RerDvyyJEbX6Ku6tOoC7ZYqMzCY4fg7RvO+8FUEUzKeys6a79L8eSo3qzxp1KlQJjXacRbt0EQU7
XBVpcoHNDfiUhbE+l0r/FLi9ZJDGm8gSqo297PhTZQaHEPVUcS4aQj7ALry8pRRKlr/WcLH5udqi
HSho4Qt3GmoFcSPV2fRaPG2DKuOs0OB9mvW0wVx9hhiJ7BYvZRdlD7Bz6+xn8MyWY3tGNGz09YSF
2zyvFBkv81zuQIm8nPTkh0Ol/T1SwClZ5F0pgnk5gW4ZBQTIxz4RRxbcskOoGbFGzgyPbGTXqSpI
4YkNGOK1cYzVVuxbqyA/5jVQFysRfVIUP0KMjnhw88oOhrkvzgfx2zlZfpcIaj2Lyjqq2OQXM4wc
v7Rq5wn2xtqgzxLSqA+nkdLXuzIcIC+YLOvj09dDA1n+ET7/Yk1gt5V1sa/K8T+dTBXxWXoppbLT
l0lNywSEneAEgXSopSY9GVJytHxongVMREC4db5nWOtH7uo8PeJ9vkAOUVB/xyQ1sgoiPNsBO8Bq
kqMGUcYycUbx4yv7ogMWldeMfnZjaE1BlYihI5NFzi61cn14+uPznAUcg2WOxUt6Z0jxcLq0INwT
YqWybJLlWRZrvmb2rF3X0INwPJLv4R/inpposKw1bs6JB1Yz7jYb6bdr6nWOk6j5L/hK+QL9Tf4T
1uGC+sV6MXH/PpZuTmC1B3PYrRSBAMfhkO/aZni84ibxUfSiJRhoauKPd3XP2xvJHcW1b28dLuFO
RVQsrLlsfEgPLnyduXowi9ob0tstIv9rSGo4lMJdSJOu/2jTaDu9bdN6RYrJ5PFt4mpfvApVZgnv
BOAfrEyK1MMFLzYjWjOKwO0BJBVrAIGiqA+0UdZppJvkm3CmyNpjp9PdJe0cJcwlSMn80h/c6tXl
0KGSqIBlP3MGGRsyzi0splg/HDJKH/ituMYg/F7f1OfA8C345bDQk+zGp5KzH/FTwv0UFL/An9ug
EW7iNFjgrhoJNgvCdp2uFbPKjnvCCfnWInlhZAAOikrn7da7b8hb8b8qCJxNtKAeWhgBGScQUxy9
WnTLdKLckIQn/F636uAAY1VlC5gLktBbp8u3JHrzdWO34xuG4kNs3xP5yQbzp4WDb/287C+T9GiY
k3J483U9KXhgokVYrJfKS9BZcjFWruScRSGIg4TfArnjGVWm6bQeyluRiGGYtAcdrxTtZD8ld8Nr
2lnHkG51j6lz5Jg7eku+W7iP7QPb1N3ovAG/EFeAcJltHhvexTJ5koZHRzBgxeX8g3ouFFzs9OQc
QQu2ZRHdvTUEnZTuc67QSRAnnIICyU6JzS2/OlSsVGFTQKtD7f2uuBtqgZH7Ium5b5WEGc6ve800
5APCbQy/AFS2bzgDj3MBCJbV+7ij7G1S86WggUwIh1znBSfgAAkrthwEzMogqn6Rvgt9ndxWtswG
eBC8LQmWkV8COGqV+F3w5+dmmOBJz58HQ/7VRMwo0rfi/CWJ/hNsFFWZg+gCkGLVD3TGUB0SnB12
/hcDULuKsVaQnFtBcj1hraf+n95D6PM4Cs+5e4wyrlw5hAPSxBrbGmJSFzLHBGfrvEuTvR1u+Tac
Z+Yb5SSxAAJE/MMksbWrSuK36FqlYP5WXt/K0C8NPcc7rXUZD1hOsTPFaTXm49GSu2QKlNrrxXlX
NTzCiBIwtyNRomwAO1pgKZJBXDXU8eaq10DNuqOcqawVghWmr3gM51v30fZLwkIll4/QXHUZ5p64
YlAOEvGqylIyvGbi7Ia1thcm1RYnuvrepyeUy/epZRQu0NYcqVIpVJjp6FMd9GWjZKwGrBFVf7w5
AjSg2gETdCOgdEk35Nij3TsTYYylIBr2uUTBBjCVsBDvMswwoyFZ3Vw8FRPNqPYmobBbixBSSH/F
NhwADyYTsq4fMYOs6aT5Fa74QE5WLdMc/dfWAyFFjfZTWM9L/fhyz/nW4j0MR8s3Ns6uHFh20YUF
MlnDX2gulgkXfOMZGp9TvTeQrUqEkgMTvDHphiakT6dwuoVbZBqyZ54OYIhr+N/H9FhYbWTl88tt
W0dluZc09XQRPsXbGyjep0RFo6c5OzHiYUW02pG94/lbb56umdNzJ03s8G+OEnFxTmJ3snEga3bp
Q54m/Ppk8/lmvI0TGVSMYmb9MN6QFLHMWjx+7lvnDhiDylMlxaMgVtsRYrH6FWQBIa0EaLOTafQu
o15J7fvPqwtZ/K7iB7j5jZdhC2F021Nh4QVY/lB9Bo5jbGgWQI2/EL1doj2zcEfBfV+mixOBPcyj
cVesjfXSQo4zQvuWTSJZWSOUVTzEL0yEjEGKQ21I5b5ymS2kTbF2qsVBB5/ZbdW9nPIJQewp61gL
nGKa7YtroSPWrMa7FF3ACE2DRP8gZFZ4wrNUuQmvL8Cx9pL58cjKTjbqEewjV8HJVNEQkAj5WqFc
x3mSVYqPN4/a7JarMVanOw7Gl7S+5IH1hWL2CGPD99hwsPT/sWQXtZOOcWgbCB53JoPQ/YqFBtHn
OXtMNG5PuZYNMnQPlqOUqLvAYoeKdoNi6LJNnFOs5V1LjQL+yANTQS/vpPeBOpxXALKZG9ydF5Uf
hqBtTRF11B1hIPWWBUPW3dKqc+C5AHuPxEJlMEUgQoVOq1WZr07l0Y/vkhlzXauBeatv26Jxet42
vVTEDXx8vjOKAgoi16YTLTQnDHro//p7F8qzGwHtZK9SZKrNdyQ+fDD9Ih1JITkBYMXK6+LfRdHx
aucMxEgfDVYhT+hBS6jJk6w56GUKYID4BahSNgVweH3BXoZnz8vb1oeD0ifgsFLQIvp3y6+NfkL3
cqXtc001GKRt+rQiTwHyNY79Y1cj6seEIzDhiWZiJuksnboF9VEdpmGEZMZswEP+YJ92C8ohI2df
9jO2fV9pNf5b/N4MrzUyG4BX0y8rXg+p4GcwbgesHpf/QUCbMT7f9DvkPBsF3dVvDbA3zhIuiMag
e2CFtNPkLk1O1bJZKrQLlndRgXgz1ScUvUbe18v6NkN/vL1PDmT1m5orkClfzkjiNNV2HfEg03q0
3L4t4qEjC8ozvzKoQEfdyCwa/Z1o2cOqtfPnsCnprFhzNtkxpRuLd7vbXUkUZJvt3vMNMnQgd8LJ
V8Edtp7EDMoWI5b/lz4skriUGNbIBbXwM/G+OZvSUevcMlHOxcgT5i/Or7RYdY1CHLdMWhKnPISC
5+s5x3oJiJs3eixzt9XnRDAajWXKPrR0VhIY25cF/HxFF67vnStZUBPnuxCdpHsiS91X6q4Nf2a9
G3rEzYYg4UuvGM3R3q8uCTsOwQH2BvLBONOclyNcJk0YHHn4BLMKAq3JzGzHbbz3RIvUu8jcAJ9a
Zb8+JQuyudXqBu+szrsrZTKJahLXbm0g7pv3Pbd3E7CfD4VXHlwDuj38RABqPHPckzQdWwgsNxou
cU6LFB04+uLEmsS+7zq30nKr+xa8c6RPeR17TRS1G3TD0Moc0g4JrBr6SxTsXL1gSFFo6mXsQNbU
B1xAQQdUvsFdg7FGtn8GlyD3zDmLBcosoYxzjH/ZBl9MvuqEDmtv8JhuyBzRM6CpGBjkn2B0R0El
sTPmPrsoyf9fCsayskoeyHiAYOsyoUnMbXaFEFv5ZrNvgXrQag3xAQ2tsOC4MNlxxkpg//tW7+Pb
1KjiJwUhiwuJXJ2FSuCCGZAdr7Erbaq0zmlhlMxUd6LnnTT3tHmkAOXIzGimhHkzYqDN4t6wVhoJ
qcR02bNzLsuwxalNi6b0zsFsLaSPEDu4wsB+ugJfC+qmm/zthQrpswKwdmduudqhcmwxxQRyS5Fo
AqYlDVgcbelhQvjAfnXRxif6jH4bSgObhKUBPWz0hotftp2/2BG3HhnxiqTui6mYIBztyXi6iDMt
UGwxwcsistDtN3tO/lkqJZBRgKqHClN028RAXVmpEGia6YpAW1XZIyElAkZCJBBpy/V9F1gNu31S
eRMwhEVKABbHxCaYxKRYMSN7T3vj37CczCZVA1RgrEO1FV62N3x8tZKXLYO9VlUjxPQQgQCOk51f
nuUDHA4bquS8Jf09HMXdSYtCD4g4CqzJMWt2UdYrl+JJHOrcstbVUmFRxSohcI+6zgvXBSOcoaZu
OgUB6RWOOIjZJ2xw2+m/13M8rtASs18XHCDCxEzCKTnpSI99hre+pTrBFxaWNdxHhzJUIpDzTo1B
TOrZP4YIKdKrdgvenNhhr5nIElrdW3vAejJcNzvr0qL+d9SncQfRoPvQGVgivS5maI1VjqrbXD9E
Xqnj+Q+RoPNOQR8kMN/uEhoGGI9LNWqQLu/xvPNuRRV8ZrDw9uWfxO8+8yAWAdbZfJ2almY34svK
nSMWRAI0tp9IpRMXBC6wA3r7KFw8dQhHuuUwGr7V63lFA+f7IXrCBZ4f7yuzNEwxUgDXEW2RtR1I
7y+oFJ8rWoXdbuy3G8a32Dgx+qUxDncKNWmqJoEU2zMRKD7CbZIUZ+5jWJdUiwc6na4zBRroGB7V
UMNncNj9d27wsU20eI3h+nX6AhQ+mv5PxBxCj5iNhjii1cPgMnlalw6MGMvGYq29I6jb7M5rcQaR
asPRKWOPnXLCXT5eHRV4paj5I117VC3a5ZYtjBEo7/RTmzkEK+9oQV8LRbSQAdud1xMRYxgBcOQs
yW6WME1QSTcEA4kT/iLy0pv/UpDiNUYe5rE26z7JdmOpi9rcYiNWc4JuqM7lWlWCIMGL+QtLYHP+
hOaNOv7d6TfhvFVBHPUohHJ9xePbHe19ojsd2ljCYRepYP7lFRlhAwvnmAfTlK5AQhNderdB+xKw
Sy2ohK3vbapq/heG6gdvnSCkE2JSfcX967SKtOSkczyQ40Pm/apCDbLMzeuNAVT5CDOb5Gody7mY
5PK6UGQW9hIuzWRPJXFxcqDUUOA8zFAZotxropHehsqfWF+VgM0aXYFW/OpuIwbuPijMbsiDUFp/
NvKC/ZOq2B9FcCvuk+PDt46ZBcDNejjBUOQ9E0ET2WHtPrnGR5ZZ7PJqxuoQe8OS7fbwlwVWuzYq
DLAcpkOGqKz/x//DqzbtH9eZzNq91J5J++/cufiAjDSJjkURodvFgSGVsnr78rCPhjGngsW3y6Vg
cRZlBXXSZISWJzWVBkq714bwA9BOQisLM9y7MXe2GNzVg3DhgrePfTscoX6lYqXN52LyVs1DD59U
Fx4hvsM2K5XpuFd9Hi2gmZDJ5q7uqU9K06iZc8h7z/C0BNhvuQDaXCm5KZES+i6833ulJJ99SQHf
o0FNGP4QI3SELwGTsMhWmC8ISp3L7K0GMwsu8bW71zlvamM9BWTJ7AHDtayqG+oiqDcRXHbeAXXq
O5KYll6MPVj6iq5PXW41QI+IeAxezbH8SMFcEGEhzMBMSRHZfy8RC89BC2x809O8rFQATg0fdU/d
terR1u4rLNhkXnrGnZtcjSlsUtWlqsP+Hg9nMq2+1HDMhJTtDKCw5RWh+l76ma85lL/jWLvio17k
i1DLjHmobZlqXE7ep035a2ss03trOrEnkMQj63AiNKjfmH3cF+JVmjiztKCU0++pxewj0tINs2H2
CKj4SlEwHpoJ3RPmIPfOYErOiMT3nVS4mOyvMDNe/xUreaBty/OWtuHDZ7Q9KnGFIdg9N1p5awAr
YmfWgiTmjRbORlvN1eCtL48k15zY2waA3ncTX4BEGssMccXw/yXm+h8LC8iy//IdtS9vPN1JZqVu
GIic+RrClS80rU/kwpjM4yiPKLhunCaFnBRr8tzNFtovQs+fo97YUEk3cfOim+D9rHC/lGn4w2wU
kYmlspFc8ygeD1+9wE5KVPedQQ5vu9OHzA19jMpHgmvwTwMPyy1DaRtKzDfvoglwH2ev+ugKdu+j
svexXCG0hHHRPLjzvzbqNSncB3D98L4z0EmY/1zvevbbO1ZVhPIMWNzhS7YoLlPKnvvyQz+CWbUr
TanAp0/WmQNEHpaIAhDVlKjVKv8xwblmKr11A8bpZwFUJKbRX4kNL9XPK0jwFAi+Dxx0kjBpYM2u
YpH5HBdeUwllKXdglAwo1N8mdmGnpaTnnbZR3EZEIRfUSaeZxzJirrQuQeJCPP/8bTy5GgWNc0TI
0EQYz0D2HNLqhWvZ+8HXk9Ticqx7Pi90vsTpkgR6ue4aiOrdb2Jml1S3uoWNr2BKAXcuY7mpf2lM
2sU0dOXsYkst9wOzlqSVclYERCj/ODbOELAP/djHDJvcqVipiy3YmvoyHBZJZtmB+0ScBTw/zalN
rkhmXJVpqdLEr8Bs14Or2uU57NIkqSAZEVHZ0Nt8iYMGTufk14Q5xkY0tocLfs+JoDGDLBwWMmKa
RfZmMlHcgdSlfyJ8nOc4UFUe56/GdKLs7wlD5HmR3RPX6HoLjrNwnJYIqTZUZGFeMw3Y2dLfkvo+
ZHeLk7zgtwj3jmqvYotgv9HrOU23TxbUqFkb75+j6wDo8n6RL+GUO1HTvolYvJC15UORUibcIew/
AhN12wTCc4MNYLzi4F0AtbLsb5Xb0joN743URzFIvTjxIuj1cb6xWcx29YFCMFwNB337dRtpeqjp
r1Cgp2VRNaWa4ILmWK0Zy1DkSBahsQwYCvOvjmZCbDHVu+a9RF4GCNnaNK38E638cyaJ1nJ0dJVt
7tN3Kh3+5yAucHwhvSwH+4AigtVYgph05YVk7yv5cG/oJnRTV4v0tPtkJDDmjLNd7KaScnYztvum
KVrKnYYJ82uEcG3gqDijpj0MH0dOPeK9rFbs83z0/itw+ELMH8yeyg7SdCviOQvbKu2mGtrEGksY
EgE3G7LC8A/1UU1dZTylFKAZNUuGjtpghsWszYYev01mqINVO8ON15VWMp0ex4/ZquhkbzEOF28n
0LtrjR2iQgGXH/UVUatIPUrL9LE935BOTYQaPu/OK8BBe5W99616mZ9czKZ8GPjKdKzf8hjGc6Vs
XDEBGt0iWXamAPhGd7oCevwCcCF+2OqEMftFCUkjrt19JuhzhIaxcN55t8Jhf7u1hJjtR+kuhK9+
hylS4e8vywQHQ5Wn9UPInja+N7UTyB9cKZAy5+YaSmKly9/oDlZe7te6n/BjvnMWgmGVR4luvtRu
j1p3XxK22DCh389K8mEDsjq0X2b5zqlOcGATfnWnAIbjdpAobYAmzV0IxXInBPR9UPuzen960te4
kz6TgxpdcbAHeL+SjOBqF7MWCWfmgd9vxMYSOCbh8gD0O9pe+wXhaFkNLWgCUlJqv3FfYu6O1qE9
4H/vZ7A7enV+MUp1Pz3LKjiYpz9h49gIXYbam43DLWvOhwWbgaGxbO4IJV7hR79ZPVp4SVV8WKyS
I2E2XcbDFLapTZGh87Kovosj2W5O+0f/qR9fFinaIvSezaKGCpS+JsCbnt2YEWLPFQijrjhBjj5h
td0JzdV6P3KG9cjirCRrzLHAeTEY4+82+rIYg3yO1mghS5UihYYH0bOq0/wEXXhEXo5nYIt7q9gY
4QUHMUEjke66ODELWzqQLmGAhSPwOmVuQrL0wdk22LP/EBt7IetIF85OswENb3jSi4dcmSdu3ooe
hVp935mLBYIsdCsZ1L9ecOFsI2EQthLkrTYpuuCa3qdHa/9cOo6Snswt1d/lAsD+m1zqxF9LPZDA
/ANSQjKBIy1EIB+RK11aYinuMhNDcEgQNpIGEeCOWWChXynmJUyROVNAnCaGpkY0UTqyMOAmXTxi
/m+amAOvi69ox8HZL6pEZsAhxmZlQfe9KtPplvpGt+91d0W1Zb1l11PyIkiaomnqADhN43+Yp/aZ
fg1UF6X8RsoDUVlNdC3K8ou2UZrFlVVKjJx+V6uA3YbeADfJJ7D15UCusNGaKF/EfkIe128/N+au
wByawrzFt/0w0mpZTe4geFqGbmFnyh6aRBVGe6e2qFtvmjwjxT5JpAeVtoVfYa1aLeEK4MB4e2n1
ovXaDxv+dTMO+wB57BpM9M3HMB9y2u4ra4mJdAD465TIrNsb5vuAkQlu9QqDF4MOljsFFHbON+y9
KMVkgbTK4+KPsr0gCYt/WKrJ/y4j6CRGOOhlmVXEmfu0NSfvjffyJTCt/8Na+5lGOwWCIt+T36Ir
oDdRWtMtqpKwFSoyuFGlwTWH9HqiGBkjjgStd/vFbyGsANe1vbpZfGW9XEnGdSo/TfJHHPchGTYP
8NKzfdbXLMJzgZmKgnVHohuQKyV919zRo405NhHrdhMVYWgiOGIltXiqxCfuhaD06V9c4A5f3Rtp
r87RMCZMxXv+ZoADA+N/g7s6a006pjs/lXWnkbdobLuzQww+YkzpGTIe2LLoXyLn5XY2FCbzqK9B
oPgtgwNkOnZYsRi7+8Zr9H6GT+th8cpiRVKuZq95QTz6QjGiE+/AUJ5feiKQ0LIqzZaUu60c9Zpy
s2iCpPcQytc+I1pffjEtVfR8454n+TZdM043dt4/waykpvWxSLSFdJNDxLZNKnhMXEawS3ZtSxXK
N/wjm8FEtjBdd0nCkx1ATohzXqAQe0hDj7u3DuH+NzvyUrZtufcIWXM+9IM1vxpBXa4N6ZV//LoZ
NIPsDnQHwWe4FkgK3BvHThe6e3P+yLLQVIzBhgKKgOOOA4nplpexqYtV4PDXaNSkdC9+OxijGJpS
QDq1b5N2B995tV9ZmJVd1SkAX9UExe28zWz9l3sEXrKxLar0TajSEYs/Gn3DqKfzH0YRWkg86iUN
CM7V/iiEi7DceVjqwR6pRMkXcMShwlJJ7kTn20UmK7dVi9eZNMTyS87SBaVTjcL4Z8E+tDVcFdcb
Q5Ui6p8ET41qcmecYlUjB6WP1Mt/0HV5oatqZvUqBNK+fenCsMvTO9DwL0hqzvgmo+E9jiCyaCtt
fMoq444Jm8TVWM+srQkcC6YYk8q2gROdFEVvDnN4yi6X7hw4t/ooHahbBfT2UzWZZCsXczkKZEkn
Qn/STkwnENrTPPWF0VveWQcUo3bXJou68a78AEfr+B43BIdAIHGrEMRGCmNKpowkPckyqar5mzmQ
OvWQ0HkeNyKAXMgYTJcNihSb1nakgAIYzo0CQAf5Qntq4ILjCU29bWp9dxvCrXLdS60HeHWdJmpd
EMrdnMRAdW5agfXKa1Yy52RfKMxichRsvdSt+h27s6iwWI+W3w9zY1d7hoinKZAzh1dQI5j7UoqU
d0Vv07VxJFQwDH4QodlZ09GtWBPCGW2VQzu0C+dX79AQzdu+yjD8eB4uBHuxJOWZwsYni/lDRsM2
B2J6qC29kr1EPj1+1AQp6U6zKtzJEtTSeLq0nZFUxfUP751adjPa7A+LSm0x/uS2jadU6OH/ecFg
g/RNuFNzUbEL/9A2U3gCEmoq4evJ22J9+vpMjMCITO744u2+FvQZY+2WUx67glTwPYctFP4Ojbgv
wCu57OsOzX+t/s0EpknluY1rCBw89ckIcaq3EGlAh828tDVAI5Loog4MpMzZVIu0vVNccaCaohNf
Np+/o+13taCpRIL7Bvs8cTf0eLyFcta2k5XcTUlraj0ZMCLImNNsOmKUDLav8YNLcMWiHefGczJ+
Z/JreiTZ6kQlIZAGLqZAmXJSE50VI5uqZJnJCMjFLXHTlFWMmpsaPTUAI/KcaIzJmPXZywLQ0fSH
i202CfIUZ0xDjVfqekWhsw35oi4SzrgpbUZJcIm9Iby3/kPAVJA1vfGIDs5B4y/pwPTgirZUxIip
3gdoQ7DDhO9e7c8sHBctZKbA3PsbR9OAUPM5JLGXkVybh/K+SEWJ0jaQNWOBlCgw4d9pbI25xwKv
WZLOU9Hlj7uwVGmS1Z9CZyVedB/2/PTVNQM3WlTTfMjZ1FLUw1A43f/9l+MWhDHznnhwZMKuDbYC
+1lKnUC5z8ojAAp/w4MqFwoFHh4rktkb+Mfff3E0Qwo822KUmjwkDwifd2KuOh3DmBKevmgi/Ika
yxVC1wNKubRA3si03vZYge0Hbd35AWFSKdMqOOAzjOXmqihHk6tlZimcs51+DIiXHaItvlxopreI
JAwXzDdfTWgMbYGA5HrP/Cj5/hyxXKt6Pq5jjDHxUzQM2R8cEyY/IeWAlxxa4LXpDI2tZco2NBe+
rJyY861Fz4eChrKeDyf7/aCW5i7I4kS4lcEFjuHbLzsphofn6epbq+4y6AJvDAS6UVgDJsT5HfCA
xMgpYVZWniRnjkLAMZZNG7Pl5V/l+cErOdCs6tcjGZHUQw/Oj/EfqcNhGr1iCbFyr0t6LJxV9ah8
02kqSGXgqIUge+aFlRlFikqb7Evm6FVP1MRgr789p3sRN3+LixX4xT9oRCW74FoNodUap4o0pYc0
MOS5BQwRjuh/eo+jDjUNHa9N2TQGGh2Cn3uExAvX1whxJF1ZZkGhEykvDYTViblaPgs/dIFkGirY
GVS/UBMO9X2lKhWVyybUsP4VGfDZHwV+RItrROViL0gWA9B1q0/VWcFpC7efrFVG3bj/nh6uH7T/
URKh36n04I01pMhSy/P+AA2AlukB1ZRtSgsGD2K4Ur5wNM7kZ9zkjm1v1jpQcJYT73EfJH/Mnxrh
g/0YDx012t87p5emrpAYYnyvS82aIZHXWKPn6y4BW0fuxnHqq3bYk4SLhQZQ4Ehr2Q86aL1WwmVT
Q2s6AJsVYptUofOKT0wqK0RI4+bx2jToZxWconKi29MR/lUNVLOU7SUcSnaoV1vyFrwnL+gF/Df/
WgbUErmHqJCkcZQ7arAWkeoQGj8DK1AyQK3lW6+RYRAY7bwuiWKG/k9cfU9WY1knmw2rlqxFqJHH
FyEXwQoPTFKuRUPZJr8o0YZipHCX9GhhYe6exH9pNkcN+6W1mtQKyjtH+nHzk1B41syCikXUZ1hB
hRsEQmzJ0c2nYPoOxaZ1khc36lYSqoEhXwqoR8hlVXExGk6dHha90xLay+73lojFqsM2qTT74N3a
Niqsy5Maaw8HwtitToBOZgUSr7kAyAw2Q9QFILv013ek5vi4acTDzX0p8/VN69OpKx5sLQ2uMAvM
u6G4Qmxe2SXeEDdFhhuhUFnAozwApHmDQmwAlqAMpOhSW7YsTKm//UWZs2o3jNRriTa99vVjcunS
59WvR5/8seWSltMMOR2+/jdGVwSnQtbjijnehikvl2BXCCVi1RAhSORIK+zTkFCkcYsX7Fv61lQ7
ZVCkDxqODzhOQj5Wm7/+1WVV1OhXuouBvAAxAqimBlF/FoP1aQOUHCes/AprJLD7vx81oQLOcDGF
x0iBnwCjFdzPWRd1yaTNI//kQvlp/VoYsFIJ08S0+MQ2FPdcG2MMCmTRae8lldYaFCRM44ZclpyW
qiQ01iNLM2xbWQpfTWdVgSdrmoyary8QkQgmts+VyYLxFIXQlPW+wxpB8AAe1jb6ZMaZhN/veAFD
oN8GerRH360ndrUNl7rI6ofV/X+RCUaKwcwh1YY4xVodJgSUCCCQ3rr4OIf2WAup6b+IKQOFWmt1
CnYKEa3fEgvIXcASrj8gIsxo5ja+ceUAqVemXvN+ceOyqAIbSdny07eYOU67BYBGpdraA/pT5X9L
xp6rO2TIAr3VyboYASILuNOMy3F4p7rbEwbbeSoSTZptGuXUimZAXiaZ1YIzo0ku8QVqiqVfTMCN
BatkcR/3wajxpLC6gASck8DT5cCqmhbg7r5wFztcSVZv8F70ypldzJVDORbfaku0b5vglXhCSa2w
eyr70o60vrRFGFexIRrroWzPUbNXOB1+ACElMgNPJRUEPVoXAl2UjSq941esxt59LnWN30PbsuSA
vgTqdF3+xzs59fLOlID66YFSOEkIAeBjYoH3Cueuk9RKAY4MpsaQcPvGTuzMQo2zLUJTX8cMnXGl
g6KCrA2VRQrH+KvaFukao2kFgLgQAy6Lg3vQrfFKo4ga2jAbUcrhGpoCK3FtCeTajgS5BdwxXWOT
HHrS3EwZZTTPa5esyvoVuldmY7kokZrt6z6XJQityhOOJA/Aee0TPsNb2nMM5GTvzTEqEHUpGxYS
X/A2VuVuvaiKjJUh8EHz24Z6lrrGnTF0+LVzyttvTdroEIR1D2a6sQmO4PFG/OD1xkGs/tiFLOBz
6XDYdB6i4xY6rd0FcilWr4BPPxFXs0xFjNokR0DDKl6KF/fBxaVJExTLBxu/e+iUCGchd3vBG+Lm
CLHIapxlBRzhQC9FE3z4YgrfV/tT+fTQnftXKLkMltg4fwceLzFbxn3vLWYZ/t4Yy+JmaxEiRMC/
uxIBehbO3OehqgEsdO2d2d+YJmz/r2ZhFZpwt1Qkdst3oA4ChWSUEn77GcTpKxeIj4dRn+HKN4NH
zWYtBNanAB4zYXygJOTXEuEu1Sfn0y0eavdCFd615e8IpBE/sZaYHCW+pNKEJsyKP2HpoV1VNh6U
GYynhd3J0YQwNnjI1vmhU4aSTNX6k3emNlvut3v/erEy7OsekbfKw0UOHcVJ96dqASqkQgaG/te+
7IAkbeE7EMfjV7wUujoQlMYosKccbHT643t0rSE2L/XVaR+W3QIjUX5YxLhmtjRHEO2qtfUVy5Qu
EKq4Dmf364eeo0962qp7by4F07RSavD+ihuHFFjpKsSLpiVabzV8bFCfQQ498D92X6jRr1SURBtG
K9isq339lpJClbLlWCRxCMJBaiAoe8uP73hTl5dfcAJiIPDVVAFO6yWVPZ3wmh7YR6/A32W790X0
qlGubRhdAKUczRr/DDsiCVe4/vC68Oy+KQ0YIcb1/yGdOmRagaWWqkb98gAOnhmxwcbdqDFaMZ3p
FHpNnDrvz4I0CT2x5AlzQaKoJEX6hM+J6Ge9Cnq25n33argHCiRTwTXuduKa7aCjtmb2l9/LuAMA
66rddz6CH9PQldEsDmGoi23KcPJejPL0/EGOHZ1Q1/nksyWVd3A/0UJH0dYYcYxa4M8ZA8Eej319
nNE57+4bxDr02ujgQfg//T5hIC2DhHFmSkYSYMFAN1X6gNOuB5ul1qt3yOxf6enTyRQ82JO/2mBA
dKVwyIc/EHBnE7NJ4TALUVh5MhUpZ8tIwrbpWicbVfwVienzpk945yiUn3Gyf+dZrIa+itn5uJFL
2Erl/X+ZhOicQZxelDM/L5q4vbHFikai2JiQtiqP10zL0qRLl6P6BPIu58yYGN4F2LFr1Re9Xu1g
xlIyff/upJCdydWSU3DiS6qXLG/g784l4v+Km8SgyqBB1H1/AIfSrB9ACRTbAXz/ISP3gA3cNCcq
ll7jGLfrNzF2plIoRy9LTzvLCcjdbIUouer77H9goK8fa/h1zAfqvN6LDsr7lnAleYaqgX/m9svH
WPf1WtABE6uSzzMY8x1ah9PU+Q1hR6MywGNezt9tr6uH7bYB6VLz7zAOFyhbWkGStiYNapR8vQ0P
xluiKkyF1IwyUNrknL0p8+BGb01dQeqOs4YD08+ifclJWVXrhNe1YOLam2irYwXMYnbQu0tCUCtk
VHeaFIi6IYh2sU+hZEVQWzyFUMRUR5Ls17sCtMG/NWECmiq64N22GdIQfpCSb0tOA8VEBDaFHXIm
udW4g86vSo8UQdfYnD0OrGRc7Dva+kf8JmE1vZGoJD1yhT//nGuifcxTvs5b/hzsooM3nsFsSms/
fM8n0bvTZ2/eNnk4Z6VNjPHGmgsOmsQ6ek29iAv3WxxKN/z/7geM9GnIWXRTLEiok4FMqVfXQvSI
kF6/7iYx8naZDcouLajqJiCvrcLeLlPJJHyU/w1DmOSWB2UUecGlF4fLCO15rfjwDc2KR2cNM9JY
apDQB3FvXyT9wkCpXGU9NsoJhxQQ1RBOGDliGOtBPcS1SQoEDV7O5MF4z2oZ1QCbPbzqfVqE2bz/
xHQqqin/OFz3YWlKvWkJHXqwHwUMgVHAX5F0OnYPngJ1ASRuR8c9Jd0E54M5dIls/+QOi3wHULY8
771aCl1aZduohK814Zscp/BPbnzBTIjhH1EDCdCZFlvUk1PtepMJyrrpew9ssVF/yyjLILsDuQNd
05Dq6NHx5b46v4Uww+dwzeMJSy5duoxWv/oZiCN+kXuVV4uBAnPUVfU8/KNLItmkFvXfgp2nB2lX
OhfChtRR9CpXBFAM0C2a/UPy3BeYmyX1KHoXvRV39Ke5wGTsAg5xo0fsW9hnTHcPmMO+CHEoJnvD
hoXQNseGIzU4hAIHfWt5zpeN8qIJQB/BD6n+zZybHN4ZeZqW8gMoWi4cvv45t/1gO1TFO+yGp3Lx
49A0C3XolOI9kBjGX/KbeNwxUgJqjigGxwdJPwKDL6kFrLUvOakaCk3fIKWCYGM//IWEHw8BwtvQ
ppEby3rZqL1egAUG4OzMaKX7xeeLXNhZaacw8HzZutd6+oPN9ZSWWhIkdAvOvAvrVGpB3kzLqjn5
v143DXaUUNdB56eoUxi5VHqGRHCUNoKrjtBZRwpyuojJlPyjhbtPN8AytHc9naPAHeaRHw1PZPr9
4lamgPb03QG+7V4z+vjwbjduXz2KyY0BW/6UM+5xTfY/5mz0AEnpvGGAI1l7KENV32IxQ7NHtO1v
FoGAtVHQ4RjrR1MOdi9zZ3CMqvRqetGVNWqQ/uxgYOzaPRtcQabNzxNd4VvFLmQcbDYckebU5Ekz
oe0amtbOQ35+USYjrVeTjHDsPc44UmW0fqyK5gpWx8p8M/z1pruNktnlKNMlnBtgnYLWM9iLS6+4
fS5C3CNrL19/yLS39hHnEUA/h/9yPylAnBiA+w4/9OhrAZkldabF35tqxWn6zCDVVb5Xf72bIkCm
2b7TyDtWd//YQM2Rg1SrIn0qPSBOD8HpJAc/FIqNuqPI1Rn/aM0WMS8TK23m1Q6/SlAOw108spjV
FVyWJAtwziA2cmY5Ugp8vKdERuBjiyjJwQLrRafd88WJzudir59oQYXEgnFlPK6vgJP2uG84oU4L
Suna8LtM59IYCG49m6DnUTtvD/XsndhovVnwtb8vcGUbIljfCpgrLqFI/Nk09wl2ybEcqzYkwL4e
jJL3lyZ4sFzF/ojmj95c6otymWkJqm/luWtW04qxavfSfA/s5a+b2TEKYaUITrYvhO+eMP9Xdsge
oTT+ZHteqOA6r4Czfn0K8hsSLUI7d3FZnLPOLMaq9DpcyaPCrToaOctVgEChzVyw+cvde3Ay0qeQ
VbWtf2O+4GPCobTWSRWQOF10ZcGTmRvs3A+uY1AQqrY35KKaD73f8/AlFoGGBCyUyrZ2J4sjQGlC
woV3n2s4/oA9W0KEnBJcqQcnlcL4TGT/ZK6NU4KCAU9cywbSs10lhbowzVtQG9TCZUJACAI069fb
bk+FEdpr5XJo8Iq9MnKUR6Li2AI9i4EUCZWcibLWe/vgXDbcGBcO6WSZFVvCt7MNMgWML22+2JHA
rJT2j91qpf4izDzvLkFC9gmd6JHldZlJAvRAnT9cB6FUAc61Vp+igrW8U6Trft0xUCLl0QTOaVdC
h6LYq6t9sbMPyXHXxGggqjc+OAOaMA1mczIxzC1inQ4YrNysSxOiBcoPzA2OL77MVk1gvdCSygK4
sEdK4I20GaYFbai2AQagQ6yslQdISF5xJB74ap+q450JcL+hoKa+B2/CnVu6hqB+GrxW0Tcg+ie1
eZ6IGoD6Hyx5ujBa4y2wFTM0usqHcSvQSenlTZz4vilXyMrYILlBzXzOtr0ERZmIz5dhhI8JGToR
ap2lqXMCobNO4bYVNo0kvOAhp4cqgjl8vnkl+5/SLawY/UDFXo5KtMMsjKzX62SBrS8qmaL9qeX5
y+5ts0ba6X4jJkFmdn9JzhMUnH9QTPG4S2IiOo0ZYRYYUjnHDk04Q6uIz+41bwDjhzL+j7FJzeQz
AyGi9ub0BYzdSRLiOqkSvS6RdjdEInTJwffKEZ8vXr7+8lvbrJx20KyVSBL5Uz4PG0NfgXBk2yY2
WpHcl30zrgVFmu62yBk9X4FDBWk0yxWJ3eSWP7uLwBxu4yvr6sUmhj22bdUknJG5aAWtKH3wQtFU
k6I4eFtFTvwL4JZFvAxbjOhu7sjN0nK7sI4UI/qlicwNxRkQ4k4IC66vsp44TFidJWGRMZpKoN/G
+kJ00g25+T4E0kpZ9Kqng2ykt+8jbX1Lsl5vsOXXf1qpSSE2L5fUbWWYRXnpNr5GhYlAQbyJSf1/
SlapoFR/TzHr2+91nrvlRf3XO6ub/dEEWMLADgBcTAmxLYJMxVJMgQtMDQ9Fha6gBcRvzN4ZXlWg
fZqyZEjry5/XeiTCmQAGJtELfjV2LUiLgzuCtChQXGNX59BvT7Vbiju9Sxdu5XrGkcS+cVxpYk+2
w2c3hZ2lrIq6BVZ1BXVAVta47wF5GFcbGaar84eAgsAgXMJkBOb6vGhlL988yVSFFHG4R3X9eZ+Q
lR0y8vqChwlH46YaysgIRuNILnHxJsrFEKm76i5jx5rjIL720CmvBvUdMo1jYfUsirOZByxHLlgn
r5dRJCqM9QzhqQQLMtYWDq2EtoYFZZI4om2c+/NmFKPV12Nvs/4gMAxFAgsn5mtcdO/GZt/yLJPE
y7o3IYNkhypRIfsb+ScZl9hEydw73daC9EM2qF6afp8AMol2rRsd01qLxR+pvOvLnEPVvNixSBw2
3a9MI/q57emfQ2m0RDz1OboQDnegN/nDKAgSLJ5YgQ9LCbzZ4FR5TpNzIzXC+TDBGXPnXArc8wFh
vwRFZPT2e9Frf0EBZrvF1pUilv3yyQd8D8qD9RHxnwz56Qe2kivnpiXP9psxzN5XqZ0pAKPTr5/T
RoTvmDE42ngiaXPgUvXJfIGGKiJbRlb6TzAUCYsIovQQzk9ctdkZuSKWbnD1M5adrDjYN/2Bsr/I
RMVivDJz62oVkuNwqAAy+9/Y3bWbCyRnqqwEurPQFLu5QFIfysVJ4pGEAddXNpWxunUYu8dosQuG
xHMCxTP1MBp+bQHjAUFDhDjWN7BgUREoVrtOkV73s3WNZg7uM8AgkHm7I3xdYzUOOX62naYwoN6g
+WdpA75ljpw0RtASdS2QblVTIuj2R1qyBYvkpXD1gJYsDFRgJNfGnS5ZZM9ak2Z22nsM0Tkno3c2
wNFb63xurnOOVDIw8QB56SSPoGV48YdTU7lbDXFxI0qu8kdBBNLKOC4KCLdLyTFt9ba0WfxYz9r5
WkKunrCOzaltUMnHcX1+UTn5NGYl5SOPWFh9XyORkjDxn8J1NYWXKSvKzoHio42vGiGeyTRhxP+f
+Pr1bSopVXwLrHCWT3JQFMOvLcfl6MRQgaxN5kHIauZ+Xm9mnw27vSevc/ElRgXDt/ZYzJhy5J2T
KX9fWJxWz2JgoiyKEffr/tDNr2Ikq4lcUbUjMYDAWxoEux1eNDG4ph+8ONaLVhc/F97kt6iwWuuD
d8OoSZBTZIagXnTbAD02P6vwNNChWqpglojqTICHXTP8smPPPmOchqK20Mi6V0aSfJMMswTeB1bJ
z8zIXo4OvXIDF/X81gADbry0ghkWgvGLEfIDX5L7JMWfeOpU+exWPTmCoghmlZX+v3U4RIYwkV/G
KFGrEYNO50X+GczmyVZrMzTDrhYSN7YMeI4VjaQb9jpl4Jb/e5BKmth73Irs/p5FhOPCimeti4RR
a6zkBZ6eXdzGXG4Noly2WtCGEAvSTEyEi+QP0ESovPSYbH+OOT0HsyWrQNNFXiFDVQ9fXuPd+W2i
zRPOwrjj7T75iZPHdmvaUQO9SQw9VeTlvuATu2975jImO0aKjKqlunD15ENKDernluxCWQ6Oj4O6
G8jDNaHil7cRhoTcohbzRKelsachcEK/RUcVRmLuC/fWI9qqtFwcM3HFJwjjguw2j35TXufpjSEI
wfstlBKsw3TeO6IpO7A72cKN7ljd8GFMTxCqOKTR7eTI9Ly68f9oPaSXTIqlWmBVUP2vVytJ5QYf
j3Ht5iX1jMZjJm9xNa/nb+3oY8bebLr9mQER0O85OVPVcMK2eGl9njRDNtazAQCJ/Wzpz2e29I1m
VaTrEs72TyOqNllCOxPdg4v8r65Xa0JvTWGP5AYXEQRYud18jAUXMZIy4SSr5E4UIZNwMdNqGIS3
2S5ogHUJ1MrzCwIrPn1TWG8SI5bxM8V33Qhy4QJlOV+hY31gvGdlKj09del6nil+dKxEw70enBmt
JZuUMO1gJm9b3G9COmByYuZiCgpI7RASSSLE4jQe8XaN3Y6cwi1NwUowroHS7eq+nEWbEG8FDPoY
lXZ6MbHQ3CtG4kacFl2TNDHom8wVrOHkB6ouz8LMnnIk6jcAz2nPmRbhbZFGtGvmfznN01Kx6qOO
A1Fl84xzF323mX54plYxig4XiUV3g9bSxHE/SExGnqW61WT/8FyUSV04vrNYbyFcOFTpQXoocy/O
1BGmesOIjgTSMka55ZFToge8d8gakPGNAyFRrlHI8HVALOFwsAmkQYL6BY0HOarRVLShOtlVcI3V
TeAspWIK3KnRWchXo1oLHjuyV+0+857xuz3o7BCXLUwHdMPD2/6f3GzF6vhxC8ABe7/4cl8WKh1k
WAAHI+8iNN6RwdCk0nwJZpFreS1zPbVqtdUDQQRnpnjPOj33rf2iC3AkGNjgnrBiCfRIV6UdLNOf
gPIKVJcQ0SYOJBfhgiUWuxPkyexykymPSy0m7BNKsEMHYCEcR5/5BIYasK360Vm84C5TZeEsjWKM
rOJ5hBFgcFkGEx/ZkSxNoVPuTb5sBsQJgIRaVX+xvkCnZ6I5v1my94Zi+dptiqRdiIQBSbS0f92c
bypxuFkptwicbY/pzfHkBFDen3hT+SzLoqijH12/Frq84B1Kns7Wvc5JspE64hltPJmb2QxkDuTS
ShPVuNZDkLa+aJJQLqYL+nOWguMAgBu73+4BgB8tifSiBacCL80JJ/9P0vtBEXtsj81YWwCBxZ32
bLsHLTjxwvlK+WRzmIOomVHKrG6WdBxF82kS6Keyajp5VQPwAIxlO824yanvBg1X8AulUs6H4UmF
C1mFu9xdTZzOwxlfuoY6gri0sz+8zNGUML64S5aC3dhR3ybL68wtrUeFlKsnszd7ok/owXsQKVzf
0bux19A5ddYhvpxy11dL1SbLW+5OooNYSQyvRkeuhbC7vbGDs1Yl8+kal6h6Rd0FFfpfcKfxFZ7F
YCDrbQ9SCqe0+ANzFoCm1xK+eQ9zQKUK7HY3NEvg/qQKmJ2/gyYCls850o8trIEKLXDwoGF1YNvf
PLotcKfO2CDnSigVNiISW9dnC9TxOlAIGaPppFevzDIjkUUXR2R4G8OXxw9ZdclxKrc5P95ftX/H
0vp/w8mKBFvVzMocSElgkmhqHkGZ4N/riOgxP/+D6NsJrrPmPdmQ7kOpNlDaOLzGZgIFfOoxTe69
y/lxw4PQAotyB5fJPlFsNaIpMSgI2FMoeEmPCcYgdRAyuL8znDsS1t9+gcEf6N4NKsaUkqznNB/m
Dt+f+DDs1w7QJIUb87b/erVOQNthiL58nxjfvRWvR8l5DVwJ36CBa1QWaYdb+UQMp/Ad++ZcF+Ly
GQR/sYgw/3/5zEe+7T1HIlmN+9zDhrfKpsnbvx/Ry0ZynvLRj4lcGlodlXxVnAtcpdxPnQF2pNKC
mLQ6HqmQ4GZwuWs68cvKKUdMr1jXMXBD4Jj4urPALCcHzuA97/jB7L7J5pmGtyZWz9ax6FhTSUne
MtyHn8c99Ly8a8/1OeSCYugEYhGjTnYsClwcKzRcRzThE5lpJVXbOH3c/wPxVsIR8ZuuJgiCvT3D
7V7KJRq+AQUc0uZ9wAgiW3QsqRV6YuPbprFjzj8BpwQwgL1z9OSg82uKpbacmLVnx4HPhZxxMa7X
t8AKcG+YYsNiBDirlwCovj7cDz0nkHtPxtyiOd8hACxDurCLo4fb3k4MqUtLNkGjqxhUoAmrOS0O
/lnB+hZOL1PPlL271CMHq4Ta81uxusA96y64EDmtmRhBKZ3Qq8Ia/LT/ov57/zZOiA3E3QmPAhyv
C3oqbaApMAS9Vj9wh3K4Px1Of0egeIg5hGu4TJtMf9PdqvfaTiQWn9ctSrPeCRCSO1Ev/c6U7yfI
oLRqf/MG3BccNw/78w/NrVPaj7Ke8qxYc+vBvodDQCz4QL5jRVWQQpv2TtjQ4f8mtszZPwG0+Lml
LXR9H/QXDV88a9Qbah0Q6yGpvHpsBFDsTweuleQtWk3HH6dliFHrv04tYn/Nz3MJjY7BvZYIQ30b
AiW0+cvwGFL6EzwIoi6SXTNardcMB+kc2OjcNuH3G0YeeGLwFXyQY6+/2IGbfYfnZG5T7CF8JyAi
dSyaEelOX3xz42b0cRFwSbvoQ6WkTSL/c7hkOZ0+NqyxxvLo92f1lPGwsIDlEyRyK5o0q64O4M7Z
v2TOstACvzs8dG8u9fzuUuV4gFQ8Gpvj2SK0ZEsfyYlyFYZM1Hw42jpgCF09W7hcIfLomgW90LMa
JD8Gpa59f7BHPMFmaG2KgvSH86TP5yD1rN4J0Qo6MbNE60W4YsOABFmZN2ZgQ9ILp5CWPiPr636q
/RVKU1iA+ZR7DARD8pxu1RJq2ZB3aaDXkvVXihfTaai0hLL+rzQDIBDavgoMjr+SszwBTgU0D/pX
DDrOccsIKeGc8R6tLWJC5AfYE28T26uAFnxLMRHS6cvDq9h7svHV20fQrlnjw122wFDWKNMol8R0
sdYnt86GY0s8wSHiyyjhCj6xtCenrRDCO6N9McRSfHMT/YleLNwONO6678Ns5vDfaT4Zz3tZuJDI
q5CEZpJNW/X63txZvOhHK10BACsMAumhFqQ6bd05G+/4pyAn4NmOgXLkVYzkoQChdsvRuiOaQ1v7
jqsxy6LambZPgp0M0wAII2dW8cjOm0NXawV20h6THhC+p9Bf1XTgj70++m1issyL6REIs6dvSoSk
Zg/FWHYUlxPDZeMn7HalU47mVlnZYsZvgvrvopSSIq3RufQ7DFr8UQJ9p++lmSWs0RUGWPpdAHfS
aZcHR05SYivMbG2TNjK/R7c9MP0bDqwhI2Wh3js1fLJzasz0ncHkeLZcuk0iB99LzaXZBVFjQS5J
oVdr9PweWfZnCcCld6YwXcHnPWJfXJO+UYqbz11sKe61fixPEsvqZeqxHaQXLgJsD5/xLPvrWsfH
l+uI5qrysnPVSBluUo3m5yXKU43cwUzrpfRjwYoG0hL1fQ42CBgBs+kvaXc4Ru5RgwYunBVlK2SR
7WkP9N4ZzzYoKTtEv+S+NISawHMvjYsyLOll6/otenR5bKI0Nfe5sOCNo4rjmutJ+2YLrhXePLc8
Ggdvn4mODS0PnXKjVVuIsfj6JklFt/VT3S8egUrjwl7vYNHoymxZVx8M4pr4fhz+7eHEJGRAWnyY
aI975APIGjlfMJbUn37m8JhEpMSRkPeTV6PpiLy6Ey1Z65sODowaOM+x3RaqY4sV/wg2CWCsYqQh
FO/zip9AGXxVY2N7uaNMMEY6NgajOMi1/0e3ce3WT28wY3uo6ilnqlP3mE1keulkqwrmBFLE4l+4
DvHgFIs7VscIe4as3vQw1oTNYv2IFKbxO0GC2aABIfYCfpA38rfMEwiE0W4NxoDdfP9JVkUzX056
m92bMRoZXI4fRy7d3jTpZYxx74nWr2PwpzcUfASyijRec2d9jRfNJWgIMuA/20hZJVNJnb8lDELp
OpVsBdMiBF2zMWffDUyGEUIH/G+rfT2hCfVgXWkCvWOdMi2+3wqAJQsKHY8xTCEVgXOXCxQAJb4+
aMshJdjEDb5Sw0k1L2APQHhvF2KCUlcFF859kRttWa2ifTVQ5QwbqcSlclWsEbOLwriuMu2aawBQ
ypX370MbBU7Kvr9jQXFbixBtj0sgFJAVICPxf7w7wEyRiFfjjoCIqTRRrkK+D/JCp+kOKsiD9jcV
9+IRtbEuGaX0bCVjWMS+t85vG1ZDHrGjVnP5X3Iw3UKimKW901XRLx6wrCsSA6DCwsLEAYpVbhtD
OWK1oaNBDHtXYelVqsMermBvBPIJTo9lQFQxP3gFQ70PkkyWEp298Yg9obWFU3vzSzWS5jRrCyzu
h5OueG93yyaENhou17uUVHHHofMajW21FbbauVwAUpBCHf2jBy+xORffTTO+SXkOM54F04LaD07k
UbyYYabpQyQAxxk/VefmKxXds+Z+jFkJ5PRoInAi3VxhL7d5v87qErVTSdcx7IA4D5UdyuqNEf4b
zp3b71yjHnM+7TusUzRTV7/0qweD0ho2O2snVfi6F2z1kxkVCfKeuvK0Ajaa1VSiy2loamQtw+L+
P4yjwLpG7RPuFK71EkpBiprGQnMVgN1lbgICrphg2yfoi68SwzK/bpdpC+qzIqXGcu9EbYO8bORO
isvXSat0UWqLwMVznnNu+BV7RkyYisI1XP2ynOGXdRwAUq5QkzsmhUWrquP58MmcvBug+tU86iLL
Dt9RYVwXxwc5bey5GZH6S7r2zd1iUZVpudcd5pbIgrYZIUH+XHTx/In7Rdn8AduOTpDxcCE9tBPb
kD05abCfpmMUfAfhbmw5Ot0IqlvodTknGEAvfe2sOY7fnpEQviyjfnFLtKl3CarkKd4/Q2l6seqv
ZN/cLAatTWwCXX8xDtqWi7iC8u6vnOcsfJ0vZekEDmPja5G9Uh7kFH/nA1H6U6XvT078agTBYC39
TcMVbu6HXflvNlXmB7AW+vTURbUVD1Z3p1AaZLU27fs5xS/iWT7Ru9UHSn+bPAPircOFaoR0pi3e
P62fEBNCXQTh1WOE+ttDRMO1bbpUhBDU2A9HeKb3aqvEvSi3l+lK/hIheIkgKLX3O3UGneTfkSc0
HmntcZO2+AAJds02nJ0xxE95lcvHzBgEHTagTPrzNXJ72kwmGTx8GBbErZt/s5xrD88JcJ+7hOhm
C/pvOO3DMX4ZN86uU2RuykVzb8zyrX1zc95LzQl+i++1W39zaktuK6pwJcZNhwxFWVIk5rr7e/0S
UZ2abwFvOSHBD+H+bp18wQGl9tqSbH+8CJUL7yQ2h0Sl0F7aQ7dECzAqJFKI8IkdHnVXG2FEbP1u
UEWSQQB9xErEPOysNRJVlrOx+YSb0suCceP+H4sB3kvJWoBBrkePnNY+YQNuBlvezRSIjiYgZkRu
+odH4P+SZ/O3pP4a7yZvTi3e6XJG3O1QpQ9wiFFVc43mfCYPWLOBi2t2Xy+tOGwborfzfo1Sv7T6
wCNqsBCrHFFC1So6MPUIgJgasmsYMYGAEbs/BXbQwCBrn6DePehdrnFFigruTCcBn4DGsdlWTPCn
Jx+TMR+uqgKWr8T1MWmSVVCxeXTP3sOVS2whA/YE6uF8uVK3RYhkgeIUFjq1jEEMJRpO0XBxkHTf
IeXxxhR3kSHXXsJiknHUvDNx/JJHr41H5PV4brrfHRaDfWnCkNRqF1E2H/mBgbByGrknqFFW59G9
Jzyqw2SCXBSxkTEma54JQAWS7x9vB5iziGmX8KQ/inV8LdNszIAv0gKFYRg9cphG8REKDEfULj1m
44QO0oYSLfkuVxK32djTAsVl4kcwRJx5U5wjZc+l8D9ZAIw/lPcTUlUtpdI8o+o1fICCVVfSnJVp
SE1mln6RPYPMHl/WgIgYk5F0vp0FuT2YoCx9u3tCm1SncRp2PmFzFzZlD/H1xO8ZFcmcB1yWa+Zg
QHPe3tRFBM/C6L2Aq6MtcKjn9PP6lknxugOon0+ENcWWtoDzSmbmtQUeWD5Rm0tDLQV9oP6GTHjz
hMrvwuI99jxcF5WpFSKD/aoWsLtNmSsQDMxxGSUl6eFvX7G1h2Cw8xWdwcvJil3KC9Wd2VssIGd1
8k60oEFBqEXpQJHXzSbBGbkWfhO6UZIsgMsLROA4CWHWe+wSb+ExYRn7viI71IcUlKQ/pqh1RwQG
A1rPZHyfxZlhDYi1uo0FAt9hQwEV8r/GxDXJQW5J68AlbjztLbf8z78NKr+YFgL90COdWpuhw8b3
BaFVAxE1eXzy0jJx/mX04svedRZD8aOrxTHuaMK/cog0OUPHdRBVUnQCnKGRcpHVVZrCbK0BXqvt
/S96HQDbMx7DNFg2skNWIcwxy3nsSaZ79StI4o4kOqWuJoa/ITBjxWjBRYEXXwi8YgxucOogzFWt
uxOuL46iyp9h8BV50FxQ7GfFWwTWon9yXxqo2rDueol61rVkyQLhzm9pk/E/5EnoAu50nwC7SBrD
SwzOoxYt7KTjjAxELy8g13PegDseCkR+FQA/MKvmGNElOGmTook7Kv9p3l0qgcmzaob8B9oECHgR
yXO+b6qN3vAZdf5yQXMV6rfR/qPmSGFLDCJOENhAGndWXidEdTOzysb4Oz+PRDHnXbQu5NQWS6VZ
ylwfodAUNL+P/FXn51eAFJjA27uOZ1FLVOVSVoRVGE3PEmGv4CIgkxTp0qb8GWGF4TrZOjfjEGHK
O3HwtdJiTV4/q8PSEBoYSZxlGOzomTs2qqYvQvB2Pfm7kQN7Y7HAj4+7ojZ44aBZrOnQIBdsdD63
XU28vKhajHy6aD3XVKjz8pJoBAgbyMNaUilKReOuYquJTgfJJnTDbgUDnXriFZmxg1kMnyIglT0j
c5Ysa8mhaoyJrQe+Kc1yv7d6OuWkvLZ+FEXbEHcBNhedp9xxv5uMYjfr2/H9yCmI5qnKTbdRsJOO
WLNg/hHju1zOU9Cm5jLxufL0exwV0Udg+1CdqDCMraIyY5vcAwH0nmVXCDzACXx5O8xbuIp+SJ5J
eG+c5wD9cDawnlhjOqF0fKyK+2WkWFiCU9R/SlzT/i6I5r4G1AlSvdH4z+q7FF2s5BUcFnPMERC3
iETMnjFLymXFamU2PrpgOd9FTYerEFk0DQKnYgglu+QuMpBbIny+OjwSTWr/Xg67tW4n2gA/Lbmd
VvgWnX/wPG2yP4+Pv4q1KvR+EG83U/oO6BMSlnDEw4ApEegNlWApfJAXCQsSej4xrHa252kpH3No
0eEqvSlWA5aMaXlvvkrCeCILcpXT4gJVCfoVz0J4YFj9Gnx2jmDBwoWnVTrHPPoV1I5dMGiJjQIg
3GM2kILny010YwfNnGL8sTXO0Ajs2QfqsH6hnjpbBJJjPPpur2ILNuDbIsmq4CY5b0GyQH6ltN52
mgOiMspq2FNt847C1ivJEmzJKcUYw6IO0MTq3mGCvt6pGFK6x8wZwmXw2QplmWHjSJ27Cp4o9t/H
I+mFRMwJd6ZII748v3VpRFNgPrHZ8Sjq+B8lPrXY6hQ5sxeOn4qn5pIK1TuSwBh/R+WGAb46WQ84
Wg9ZP24AdaSKlyB0TzZrM5XFKHwJvfuMTWSdhR80du3hmJhjlvGgd+CyBPWRKdx8oi2TGlxIXkEk
Zu8CH4KXHo+PloXMY6FkaYm3SG7QSuh/Pq6LL//cdAmQiVjxCfYEmguSghglCIxzdEP1YBfVLn8W
1AG5g0O5xT3WupFlLorCzsSsT7jx6npZS4SIaWOJi+ghE9ftB1RpVACHVOou9Llym6zyIFNYW+OX
IKgpiSavDvOWApsYtUc1+ZjzxloWz/D/W98mWZa+Zepy8QXgYtjqDXWAMVqKRYk1WW8XMVF91B+h
AEQ+6Gf570Kqu2zMMrKu4QyUIVZ5OwLyzkJnP7tNN5bqvMbIlIbLKvlkUYsBgVCwB/2ZbHa4kPSQ
NEu8wWQHTzPYaVIzwS9knXKDC1nOX5ECYeV5ExBeSVd2yqh6D/YJj6OQy0xsgYC8U1UPK0YHzqZn
TsM/tnm54qgvtIMfrn6Px33TbTSOjjXnf/XZ8P/CYbBYCtLFIUv+pRBUsa1U13tnZWA/WlT6toSS
BmF5FBBOiI35zt4Jkd0JwkKIr4lq3H2qmEw8iRp2+CA2tqC/GhCYR0CRqk6iWyzKDUSWXZEsG1RJ
w6o56aS44UaD5rWAGDchjdeZmHmSP8iLpAWnSxWB2uzMH0i6sWP30otmRLdj4En6FoX9lFKKD8pP
CCvry9fO3uZTfyJwZXIofSwJTyClRxiuGK1mnqo6JrqfxouExrH7tr62CDnbCAbh1Sy1FQDrMmKH
De5yWWRZXojsKk3b/GpIQB55AP202wZBDTlgJP5U2HOc9UIRxR6vjO4euyKw5f86lmXPK0SkJjMU
KC3b1v6WzfHkTFXWCIBIODuDEx7xoC9d5niP/+ROTvEuq3WiESONvT8LzQfa0KBLw+2vdYm/HhPo
eBc6e1y3N8fZjWorKExpXCM9m30l3MJ4Wweuk6OL/9viaJ+yRcUqhIZ6nxxQUIen+poZf3xXXa38
aD8BwfLhu/RrZJ/AYGYWqXck3oNzGGFMbFskYXhazJdUs6D0sKAnjzn6E0YbFbnh29cdkMKbuN8Y
9680t5xZdTP/vsHnSTVcPOXiKaz/j1FgTfPP+F59MnTgL7zUwyvnKUrDr8kZP78ADVGSCVAXfi6U
7d7wR85U/YTp2KPdd0BHzsMhDGPLNWXgBl1SsTIl1EI3HvNLbOWK+b1XKRXD5Y7zIGExShJzg0+F
D/FtSv/+4tHSG4moZLM/uprMUqENG5BFa6/IdIk9Z/W84ckDQSRMMB7FXFczFEu+tN/M2tkOdYIb
czXpK1amEjq+Fy1LLN9SXIZfNPn99T6qTi0B56Qk8i69fSsKMmYsu8gJ1zN7F+Cu2EzgGq0El59r
dF6x2CP5PAeb4cXlxbYxD++9pjKpF2M1smi+bXZVy0WMvcZaowsRbyg0teQHzhYYWej22Hzr70pK
7qSr1pMyUBFtkdn14ba12/xiLDaTOdtRcwIpJAgzzgsaHFRgu2p9Ht7z21T220AxdAG0OprLjcJt
pWN7Y3QDqPHiLWWm6SD8keEP5jNyXtH7daUHS7RbbtbmrzkP6DC2Dy/2fvc++qySRvY9J9F2Kh6Q
xLNOINnAFVlU48hU+FhAb1IEKDEvB75sb0A6nGfD2CR5GXVpu5CIdvJTEOZNIrebVRQia+cuxqzq
nbAKdstBTsLvyTzbppuM//62bASdy34+J13RVY7UaFkkNfWrN/cnZvw72IfYgHIv45AlkgGeTl9i
Q27odVEc0bTIVb6q/vqI5E+zn41nicFq4DqDh4Iqh8gNnQ4eHdd4cVunf68WR2j1ZqIQF81LpYC7
fkfdlNBYRW3rCIIxYNhh3iDXsm7jbsE5Jx652q+HzElriPCdPSA8teXEBoYXtN+NRIaPfSJj0pg5
2q2zZiH4lJAhF/5iwG+DWzp493/fiiHTXxzfh9vvz47aqoAtedjJZAr6l9oL13BzNVCFloSsq9Zu
G9UF47W7+bdBqLDm6nuDhhvAhTRDABdx34EfPIO1KRqDlball9D1cBVU1+8I8AjuDfAfax/wAATh
o4i1iG4IAJGxlLDJeBU6SxM3xd56httbSa8aTJvsAJ2GHEWVkoLxLKsYrzsXZ4AzQm4blUCdqFA7
BG8uwmCY117Vn5HxdyUjwp/qlpQhOptP/48+KukzKCMXp02GWpxGHUWxTQJ1vNhGIua2us9i7erf
ZQ0o08oqQ7HD3iQ9u7C84XFgjgi8if3ntkzw3NLyFKPkD+ukXyXyjMj6lGpqydJkmIU9c85D5IAt
V1IMfmN9UK2Ur4e+2QjIZwXR2+50+0n49PlEpZVPtsNeriO0VRg3BNeqVhx82LUy1T+lcTdW/DRt
S62t1YMzEvj5IzqYRNH+h0zB9+RH3kIHUglRmdwlH7ZAxyY7XRoQaXqA63MsdbdTIrV+JPomkfY/
ZDvUWFGW9ZXFsEMfLb1YAVjGaPxBRWBYhO7Pq6hGu8kHdKxw7jlFuDtmzdQyQJ7ytz6UaotaVSEu
5FVHuCXWOCgzh9gDd5NcOK5XhbKmh1LAwq+s4fu+ucZManZGVsxt23M5CHc+XYoz9L5DZQLpM5c6
HsLJA5Q4AhRzIjC+27N7Bmnx/N/qP5yRCda9tHm7HgGgKnauDqBfuAyLgzwt/6MNcQtU/JfxUw98
RFrnRoztlFCSucINuM8OOo0bBux1s1UvV8sLcUE1YkZ3SVBPZzP+nQNgJCCdvs8Wr2LCIbX6Lr2l
e3slkq9O3e4wSj+yIwFVkN5bS4a4C8Mp6k+EeVzNn/ObtQGqepvSj7bU1EYHUNPOXb8nu9Df8KBA
yM44fJnetq1M4btCrCDGAOZCDDaRAi6+pU+Jt8UA74xWhPGdF3R4u12B3NCPzwwXElW5p10L11iG
XvlJC2uTzQz4eIPeG2/PFEulQZPRBukQLx4887GTLYAuLpv/b8j0pEHK1eel3AYFLIEQ58VipC2M
7cPrtYLGLMXhzM2IUxC13D//XBPLhBqO8VauJayMT27M63qzT0iHpLwhQDnwCRvBS+9LfDDm2Ncg
Un9EH8ooqv0KZZwvSs1e0ru9WnDBXZ9+Sd2rXzFhUt97yIxw4bOneSYmAu/FoK7fJ6Iesg/GpPYK
pA8dHEi+Ugh1cPWsGt+DVY15Bq1oZYrzOD7RpIYgnZPLBY6t0h8TPMqtF9LvfaF0/UW2bWjJBM2F
qE/SibeOmHUw58AYqgdQTpm3blq0tCkJf84fckrtt1ryXw2DlTnstFsAgRMx2+ZD+8ISeTRJqivM
FirWauVZ0MSTdbfDonxTwT3N+w2Ojy3wAk6HJAzosD+ZIbNrPdu1YFadxnm6RDzuUZBFWyZDZPEJ
rGCEzuBgAyWavm5LUEniizKJUuq74XvkK0VmAN2RaWxOdL9h/SAVg8yqhaFABN3PdtLq33pRF4jB
YNgaBc2Y+LLA7UKGWpavdkJfOyos/M4lrtBVJCGuLwwY7x6i3CRLNqPTgpewSINZn1bQYogz3H1X
ruNvVi5WKXOxPDu0/KqpXg/C+30nmcxsfD7CjxjVv8JR7+2H6rDXDsjUlhffAvYCi6iXLkcPlbaO
+ggBmua+WNCTVxrd0eTIhspRuoIedIc4/aTDUDvZBOl+crUDYGuRxO9CXS1/dGEt/TEBrVL3nR4K
fq2gmXScfDets6C7ADY/G/zR385YAGjr8NiGJHtgokL87rxRdlv8DYGnCXNY588O/f1KyAA7RVyW
mMC/8E4RXKXiRgCRg/XXuDtabcE98MQz082QlLlhgggk9wUg5XtZTUeOjcZgcPGJPU9uJzdtG8dl
r8Ec/gLW9TIhH9Z7TgWvU/5nlLvK7dViMupROoYhwx/wlwL2JqHa5vzPdjSwnAMvFmqbJPnC6wuT
Yx3z6ktPWFnt8M5+/0nGdiwf3Q0TNUjKqV0GMYiAhD0RlzNhUu1JSSGdm8TiHq9KlNvI3pTUw5Rx
9CA8UUK+bLIfqsXDG9frMP/pEI3dP9/5rCLz7OOSZA8dRRaf4YdEkrXzwUmdWJvCbuHN/2HgSFUr
wWyYivzEshrH+bQIaKOj/tnAbitr7arqGvGStYhSUbxCV7Ir0jy4Q/BRqOne4xR8+ecrkx+W5FCN
QPDTdQDoqJ4b90nOCsBk3lcsWJJvBAn6SAPd/uYweglLd0Q82EKg5oMytGWmVKK7w0XPCc7W9VD2
nsIkeIuT+6fwFTeStZQ5lMRjkPUMELM3Q9Z7jPfoA1szA1unQzv+aLa0W0AqjQvSp0HKuKgeuAvr
v9gdSjGKBoarOECv4DBk8M8I3uDd6MPwDblBAXrG/hL5BYlGA9XTwah63A91Ra2jgljRUVspHe4g
JNi4B8Snm0rDYYJg0Eec5SJeYxZOX7VK4Qhl5mpyEe+vLppfnCnoTQRpPbaIH9gr5aW+eMiB8kaN
NYzxPrG1acG7pCO5OlnshE+zgSuXq16JGvLTEIbOZQsnhNgB7L3uON/fSxEiC4M6jCfhCFWEp2GB
Q41fFm6N+zj/5Cp187bUw06LvEPNP17GgoLHJ8/u825MJoyiOsCBOLrWhIgkKs96sO5fuYtbLJ7i
SB1CKyndaX0MhYFiwEi4geuVqah7hax2VcTSM/BtA0FwQJA8xXwZq6S6ajxwAI6GZ7PEwqhcgU2k
tCGb48gax7F1vH6lXuQ4MylIhlLEZJXC6nUILH6Dnk9Lh9I4YOsTErBknren8BFnkf/bdy02mq5P
onklSISw7Y9OKuy25tgUjzfx9+/lc8RHTd0vz0ewN7nTn2l5cPuLasWpUOwQ/ZH6bT5bVDJCZ1R9
DwKPDxUQOxJQSvLkyfPIL4Az/Oq5vtvshPPFBxyLZJ5ltPapXmaihpmXarDMLNSwg2UqTwbE8nXG
8YTCmt6tT+auvDbTyk5K+Fzssj9RLyDjh9SiQSVmR1+H7Y9+DRttJQlCqeQfXN5V2QWlcMG+r7mv
XU3g62+GG9eQP727C0RoeqjDI/gXT0tosaXRgLhigYzH61cnUDCh3Pcp5muZEy/YiHhYpMH7aMNH
x6AIbIRBg1eXQ+tFdMAf4RUTLqN3WYPEwVomLGeD9Q4G/i3AYSe3h6krQxkrs41lwTNGocYzH2zK
jrR+Osbx20xfM4FqwaZUf+0quG2wmOXIz168ne5K7bU76nAMQ+TyaiLGN154XE44h2/K5ZWRkLCa
bkgoEanEUTdO8CY0DJ5As56Jp6g4KkUjSLCoqX8iYosh7vNCpLP3FCsb+/RJ0XFMnmO5tujHocLN
Z4GKk6v0RR/f/ELRd2q3jZB5acg+M8WMuYAUqZOB9qD8XyBtNdRlX9fUkqSRzC87Qd+UFGi+q318
5+HijlqQRSLzPhd0+PIZHZq7c4RqCXYNBsAhzovN4xFm6bGeQiTOKYr4V5L2AdJoevCQgxPjx9Bc
DZHdxVtBJ1NKLkUcrotEvG9dXD95ZHh2Q6xM+cwvfQH3f6Z5T/MrKpgtRYKgH0tfTMZp+yfDYE+S
4pRx1qFaMKDu+UdbpP6NOpAZ8RCkO4bKJBG92zimgEgCBdbeXrPxgvkoZzO6tlG3N+im+qfYHRfy
57EDJLaQ6AUVcNlfQvVebvsi7JF03CnyYxH0in7wsDq5/bSxZ86qh7jY5WQ/pS2A1EZEnxgMP8/b
0Yc8K7O5+5yFQ4bwYSguFB+h7Alg+a7NVeHtwKuQ/f5qFB3Aqgs/BQtX1hrq655T/ImZFfgLskmH
GC7XtLqEqlJsZHacsOXcu4l58ZELfqgPo2EVD+4bG0vKg4zAcmVENl+ZGqB4VZiYWYBFtUta5Tzs
s22CArnG5Z00bQdeSbHfR72zEn3VxV+zoYD5uAZSAJoHN87+2kqhUL+9c0FY93jcfKPPWhtJV+Ew
QgJsVZi7YPlhdAJX5f9F5jvcH1EuxE1SUp+CC5HPxgi3qfU5f9vBfTg0/Hswvp/3BYNU9ZxAcMrJ
Rn/7K8vml6D4D56lcfu9iFdYiM+ATtMgfL4vjkcY9IY0O3EOseKSK+KXXUgCWxi1FaNMI1VI+zAf
k67lBmUMLfp0n/7oDSCOizYASs4gzJZpiKsujAhi5HJRuG3NN/mc3hTlTIeOwLyf6noWGjmqz/OE
jGKibcKiWG0joyUgkp2axlA/r8KZHGMyuzIQY4tY9mzRrZbjZBLCL8aEigdo6fAMcGSjhS0hMHRX
NIdRLKjO4hqHahGfn6qAml3JKtjNbjQhgJrpjgc7f3VRSUQOsqAXgp5YqchqbOwBLDe7K8Q1ebsQ
88gGCZ6Ya+rlKDaHoc1DSZVyNJaNAFHLYzkvn2pmsfLH9u5wPO9YXp8IbWDyNDIV1fbctR4JYPno
xXpIKs4GjdNYYrHYkkT9Nys9JP5S9XbgS3d/KyijXLoEHbx2NseKztfTLM+9ABNEeLWL8aOU/qXw
GRVgvL35dReBdZnpOG3+Tkr9isWnwMO6SIV+yOR1MHEpP5lXCKsKYlOLOvo79K5s9sQdk9xS0yA6
FaEk/loSqZc29Cd4rc1TYgmjoGneFpGts+Fsn9FI8F6ppHEuhMiLEHodwicuDmg7vz1CK98mKLlg
/aM7cqrookJz7mHXzehqKzJrTDhxGq7n2aivZ0nZ4p/qEFjT3ZrrEt/AX36BjGFkCJN5dve3MpSJ
IY7tj3rQLcY8Gqb241OzFMwDG27t0Q7+ihNLBnS5ao5SFtWhzS9pleY+PQP9gkBLpjdNkNNLSCVS
45s2iL/EPCi8UQWsF+Q3GGSGnlKEv+GK3QzHu4yIT1SEgznJQcIzveOCJo6Op84yek508Q0ezsqj
UpQAgfb8DgMwDBkTTVeYazG5dd9eIMGQszSSdJDFYD+E8X4iSiX2m2rm4C3O/wUQyyUYk7xXk5LA
wzOmxpNDmfGHGDVWCUeti6akxRF2k9iAtoF6D9ddkBU2+2wihg0mBXtqCKGi4t3+YrH/v32/uO3r
RF0/EEtRR7btgiMRr5JCWbxkjAEJwIMO2vgLIT/ekdrWdNXRGNIBQPlA9L1tSrT49DNWIhNbBLYe
JD5xIVPM61Dwd6qY8ZWr+XvRqsQniGhAaBqmfNJZH46cTkOq/sTDESieMBY2s1pVaStA69UwM9fl
uqKDbiXXwED9rHyu+EFkNQXUXZMDEizqp+b6XGmISo6zadnVt93CzLL8xQpr2CdTyS84BrE1O4lu
+RKoR5pnFi4OLHXcIo2tqUSY7lzZovPTTn+a1kUIC66yFcJ6iVamv21gTFFid9hegxZSeFTGnI+q
pRVRkrqM81FH7Th7YxwJeaGlfzI69jatczrMsO+k54iwcNqzjozOrEMlXuY+BhujVlhiR5oIsMhQ
XSV1HNO0Q+uh+Nmtp3ANr2oeDjnpeIgggH+GTlwg1Yck26iRLFpT0nXOyQ8goNeuk2X3kycW0gc8
ZP+Hz34rEqLuOYtt82QRfiQQfO2aXOBGe+JPhO7XNmHku4dOhOzX/5umpre53QifxvpnLwqIsS+t
Z//YT+Apkr7KhI8gsyOsY8TWf+Usy+LViq3HFoBLVhsDenA34PqXBctAG9DlSsvFOlgQ0qVauQ8v
kHg71XDxXL3oXCRPyYnOMjRGqWD38yeNV2y1aZ7zrIH8vHqugJZCNzUilD7kDssr8sgc6pDDFBN9
3lKT5w/yJCox7uDKmNQM5jLketILy7zNKlC07HZeQ73HMFLU9+efgIgLtnzHaTOY8w0dj6gCH8pk
aKH4woAHmElIZLZjGjIH5hIsCsHBkYV0i4oIRORMGLHR4O5IjzZrlRv58X4uPeaULxuVyhBiGFDc
k+6uG+Jwq7+7uRe0AMpfICSkp2d14/pJEx9zgHk64nnQMvBuWXaURRniN582x6gdhmnHTGWyXg69
PA1gqmT4EFGHLQpbXs7sLZjc87Y9Mnhwdo4Z5QNL8P3xkV1jr2EJiytxOtxjrFiG6FzNy1OLHf79
EdMOA6aVnUUcaHDkiKP9Vs3BHvvpHKkbd8xgh6C2sUjXCmSFT6qfUrspqDyyb2burwVN2mn+FvOc
xU4KMZL4SXGeIHxXyQrJwJ0UKL9hOSdVMOOKI/1uOppqOZKtah/hOwXSlRuNwkhVmhND+c31Rk+Y
GwYTTlQqYwJvVxBDO5fN7QGhNTl82JpouiLBZQIS7pbB/jsBsU+rtF97DsD0ghX4xSz9AiS1+Krk
LYxD5nhQTFnfKe6IY0YzsiTP3wSY5Dxu5btUeQKUqB51m3vGeNaoUCb5f7J5nRLSKIvrget1eB8K
jO5qy4htu2BXYqlQFOTlsjvFS7vO2ILu8SIMJQbjFwq9v8Canm5+q1cjv+SgF1FXAhQWUFNza70H
Vl6ngCYsKmsfULnEh09EB3O0fthPIEpvmT60ztjFl/bsFphhMycw+RFinMfvfOo78LXS3NFzKhbc
zvIliqVQ3PmXyUS+QEQQwqdt6T38uTeh6H5TCZBZ6F8Gav1JSAQxgcBltKNowv0la156MLrFBGsl
wPQCXed2Ey8aN/T8CB9kPjE4HX/Wzm66phDf5aT0IUNs/vLT69atxCAY77Ho2tGNqNYsJ8we6M29
7hrJXGe7c7QoTRt2PI5FnKO4HTercXI1+KDBlzDRIz2G4osoe+bXgwBCaD3DxT89y0m5FWs7CBMZ
fI04rNWSwWTnAuvXT0BV9iyw4WPfcY3jtg6gvl3HywtfwiawlwS5jj33A3CZhSoE2K22T8Y+TupM
UFkd7MkgDSsHmL9jJQ+NvYnw3S+XJKAVbRTcEH496NxM0uKos6A34uH5KY9tAQmAZD4wM4BLwv3C
OgSbCYd/HPfJF7fbHvJ7Txz2yKAhDmbGG7PJcUMOMRFDBzoO2MMi1OMVv648e0mwBpRdOuST0IsS
hKUPgOS0MhwJH0barQL3hkdwyL9Q97dlEz/ZumZv9L5kFOP5xQJYXeCIgAvuGarbFQfQSrCrUs1a
FIwCQG/0TxKuLq9rSfIeKAwzRKzhp+k+cHGT7FsLGWoYMECqtZtExKqwyzJUI0fLWVVVTzYkDv/3
x2gq4dTXLZK7nPYpHEg179KtLHGE5/TzeerpICdMgrX+JinE8fMZ0EVHtDq/4l0tqMpVyCqpNk0H
XfzBIrdmbqESn9bG/BiVA3bIwwbHsSm8/04EslF25SeTj+VUx7LBzR53BexG1dSffKsmXRSp6eN8
CIQ/6ihTPFreJ8o///8euR2nY2taYzauWvLawVIfg+dMgO3M2ZQxMfBNhyfkYSVUmBSYl8H8LIFv
xR4DvcpQ7bmba4U3huvz7r1m5A7RAPxiT6hL34Ukt8uxzVllAQaU6tCLB/oTpRsDZNJLMqWwMx1j
GO6bZH0m9kjaVBbmgOMVGjRnQsAlXMaFASqOgKiGquOo9N+IzJoil0KJbcz7oV4PPtpRuKXvkQiE
W3N3HmKs168THAEBOPlWMk1zkPs3h6nxtiTk9TD+kS+6RLS9J2BMY0cEkDBKcmuiTMirXDJq/in+
xsQaH8iNZ4AWNolJe1G++xF9gChZXKhyFEbsJUYVkS6pvgYETYvkn9NGHoKNv4h6Gr2MYv5hQhUh
/MtxNG2xbqRhVZmOWTntYH7UlIOpYqubLCrC/3aHfK3ZHOx3O6rbcLuhdN4qNZvSI4lV0rJLHxN7
otWnuM8jTAq72P+tIenzlesVdQNAH6K4VHxk3hOv5uC0p2/VhRhyNf2U+cDpiBBQ2IEA8fklBUGE
oc2uVifzYH9EACzlNu+5xvhMb3vpVwdLG6iKzeXjZ1anHJME9k57o8gErc3QvYIbrla4BrzCIKVO
K0HEmwUjYagENaoInw7HARLDmxhb2sz2XiaCaDiZ5losKlZ8B++qOARtgmkq1GdIz+05Q/yV9sXd
Fc3Wo8JfZG9PHel6tkYktKB6cM0mfnnn0FrPgq2EFsE2v/yS2WKVvplk1vkh9DfGO3WJjNQipB+1
Kx07E0jGSJKD67DXQ7J3/kpQRv5PLcnD1ilLITeYNTyr5ACH2d/RIGe6EtCmYu4Uw3encH89F6Mg
JKlmqhrjAL6cZpbmnqrYuTOc8/55udiN3N6X7k5dABk+/yCnNAXpqE/lhOdAyYMMXd6TjSBhRAiu
vj0M9j1zMXl3+yhuUeybeusSWg0SYCx4u8sLz92waGM/I+kyUbaQquzsnExLdMeZJJd/GkMJg2B6
VuFU3gQZqUa0h1fyNjcVtc+qCl3ukhg9YPVlhZ5P1zOkh8GersWT/azzQBbkd4376RUPX0m0/sh9
5eiKjOGlA04xTSG8zpuDxkEkYhtX5Unewby532zw6pwN95Dj47QF52BSdLmxIw7qnXlqlIXhG9cU
QDrDoHKTVMeTmZlk9CMui2KszUjo5MqQeoti+Xl8LYGydUSKYD8H+fGfeWrkj1gH+PamKDDl9Mx2
MgN/iLE/Sp3blrsoVDDjo1Nsg7LYDyon+SDFhHcvsh1uc1roDv7qvdyCH0Mjk1/NF0NCGRnIeyre
0pPiCuE2aTAvgd1X+Eu1wZjDd4optp97I/jkxG32CLUGah617BvhT26XK2xi9IGE+fH2UmIfxEUb
fFq4eaum4ol/Xkv8yWZ6ESuQZvp7mXKRA4xzZth1yEfePs1TizMSVUGi49Dm2BJRnMwJIOEe1KsE
G234/RgEKABMHLQY4TOqzVGKvWb5oRy92rG5Hdg8EJ0h6Fa0kafldfSTqfmSQKsP84QLaVIe2scu
c90jUrp0fyji9Q+NVhSuWZS5pCrjSb/U2ei5cz4U3hK4pIuzTGrgQv8b/FwVjth1hlByF2HQe9wr
5AMVgNFrUIyga3gf5uZZ0i2EC9iZBzyj0o0fYGmGKt4XcY39hKD+9JkSViy3yZODJAP9CW6iWCWQ
ieU0ieV6wtnSTDVyWWqPxvyOlJrygRHi/mxi1J0lohhUkq/qbCiCXnBoKsxI96YOsdS8ZGRwbT9a
IKhqWZjDdjzQWwU0n70PVb3rlUdHf2l+5umYxW9k/C0aRdN+ech1CoFByNLCCEbIi/mmKvvOsQBM
FH8qo0QhMXNHip5nAMoU8tpnopJ+ym8YTiHiPzcH5KElwveVIjQhmjyCfO4SjR2Yt+E0VfR+BkmF
59Ile8DdpQ1n/PXEJyUiyClytOJ/R6INclQb/tFpX3tk3TFtQQLKc4qtJIddfqMYarKrug7HXX6x
calRTiCv7KG54aGLA0srLwu1yjLFslfF9nVzs/Nfsd9Tpr1LCwnX4EVk2inncQL3D/18SEhwEbuD
QEdGE7g2RYCeeV+xOfszbAdsG932E6512aXFWOFaJcmzxnajrCprhPZjgbZKqinO37WC6KBI/HxB
ObM8VkeiE9TA93LLxtuJUD4P8mSjw0DTOa1xDhLVn/8lowunKTkRhcKKJv7L/5pIp74PhyiD9IWh
/8/n6yR1mys00+TUoJeO3rFuNr/r0r97WEvnAv7HNxPMzeV3/w6L6lLQ/yfjxxsVLsAL35Y/8U8A
MnvW1uazfbAWK7h53NVGfhrMBPTJNTE4MQaL9LEQ+RldtQg45L58VxXGnH61FFnt2R0ARmNgzOCH
aok2txourKKzi48RUCuVBjf4mYOq2n+/kOSL56FGR7I8lLg/lxneRXVMlikKEmZf6pKR4f2FI5E8
tmRtl09/Zdr5Cfi3o5RLdHeRGjnit7ne6Dasr5CjFzcTxt1JXBDK4NB3QltGNMxPNtnU5KJXCyXs
t/1TjiGYHR36iEIEIj7DMYXKvH5Fc3/NnvVn85OPQOCh3/TMAzrsWI+5i3K7//Kx+5p2Hn42L8iR
tSXWmwP+RFSBUPdjflccLmv+X6G5MB1rfR2eKfsdQ46en/ir2Ty2t9amNUNYiR5zN0yHcL+isbmX
yLL2LiYw0Zv4fycqknoNqD8cjSTsaxAjauQ2FYw0TJMFXuoXkfQTye3j/UJKphy1AbuzygfRNs9i
C1wC+sFzO3eG8FrVXg66rAB2bgdhuKvpiSfp02lPLC/sGBDX864goSXHKNiPbrzpNPTrFWxBtykx
22Z8h4UXBalmmUEie/suhtWzrpjkx7Mkma+fcx/04u6K7GQPGATaSIjoXqBoUlx6ngBs1Z5h+kjZ
tn2FoaUHq8BuVWx0ws5L164JGboE1hptk7RnGcQ/uXC0uj2XwaHLl6IyeLLuriCOIDvwrU5GsyUZ
IwR8+7WfoJgipQQ7ayuGP65k8Ysw/asc0R2k48xI8Z5W4wRCHIWvMYm0U16+GryQiHFSuf5I0YNc
uENQJBOsBc43n1yw064bpZyTE/vlO05p0V8w39wNHzU3KyeREwstLfctYXLgFMMRXNo7k35r7Bto
QWIzS8J9/taBMaF6iR+IuT7J3cSE08tdoHt8N6HAyvIQBLupPKtHzu0KRI8Ne8NG3hsLaeL0Ys+l
UQ66uXONm2ZOqJBDvRL8FRAeaLfpJ7MwQo9AHAAqMiHhZ1FAesX/t7mz4pJwU57+fiPLLFu00Enc
pgtbmVJr5BLwPhtdHrg1Nsc2kXnfASKrKjgKyDvzujBWAzf0AiWYxyEx/SCMRqTI2CUH/mHx4mSW
HX/U2LRXYJJpU5DZaU0RfDWXNZRPljLIFHDBPKhUBDmDSJyQi4+iRQZJodpKaJEGvPZx0etxuERq
E8V9Q6otR/VVFmc+1GmVRi9ipGOh7+tuxZU8s+Ja1jRztpoSuCv+Lk33BPhVUiCdjbW8OiUrSjYU
/498+NW9q1yPVJrrauPLjK2itIfRtkC85NxSUziq4ohg7aAu8Er8vvYlZyQdy77dwpwz+DX/43vw
8HYO//MYjQjR9XDWmzK3pkMnHtSqEyM8l0MljmOZbziuBDkpycW8z0QstXqh7MdduYYBtNa7HAig
7YvO9clIwPGI4jDXTUDJ99Kx8HNMZrys6g3TIGiaE7eRtdR1Mp3kLdLr9cNuubmEnf24bNWOYvai
jT8mtn9ik+nd+8l5lV7fEGMedMcdYXdkfZHxx4boFsEYX/KQILlInb1D45cNubz7jdjHRT9NUZR3
981Q/BxqGAzBh0NvHqPse2sGu4BWw+2QV2hhcOemSZDeOlLgbKYRo3Z6gKjpizeRkkvs55BfMaYN
4lbiwZmQHDlIGEdgMKTc8H6v6B9KQ0ro75FWsySWzfTGhqZs66h2bzplYQbyJeD8cDEAxo6dB7ic
KkhsEDF433sMM62MYqYmgZ3lcMzf42lClDd4jfWF8sC8372j2D1eRzMzjvHkMte6o2c5MFwKFdA5
jQm2Tyy/GTtoVcnSsaHFFh82ugsBfZfbH1xGkSOoZe5eKQ49b///R1+PTKveuHQFecXcXNabEt9c
krMthHRzu0QlsDxRBoUVoY/g44Y3m8MOmBmC0cP/EgDO/PJD/BuFgT3sGUou66Kr+6iQl9BBwBMf
5FYiDtjUUDYEjUK3w7VulZJJmIzDlCDV8vLzGTEg/Jred58wPXTz143KbKMx2Au3hmfyjUfGfF69
BDMjBCW04wuQODk9zQmIpG6uJw2D3vph6dLy3/I3vDRfG+i3tuItN+d75p4YGGiFL/czAeoeVcbF
Kcuw46vu1jM67FvNuuV5UbPPLqrBigJ79Nk3a0yw0a7JHb4ZfnjQ3GMXL9hCmrc2Va04a61SbZ4g
6sWMdNTYiNli2ZrjNGIm0HNMm308ObVv0cI+rIynoIrgFkDts6IGEOHLyyFUyoj1EAGtY+8EmFMp
JB4iOPf4QTjI95J/HudnPrjPhitVUem6DGn3q719wSVAYhcvU5WJRL4uXs0byIHqEB2AQpuYfBjM
QHFnl2mMFJuZpqpjSQ3+xJlm+0yEKpjCaIFHZdLPKIJJHRxih6zZ4lxKTD4D+DCF8Q0RY7yzjrDI
XVDXh8A0GxH45RmSzyT2EOL5MZdP9vI/Hjz3e9js3SR/VPla7BhTYX5Xi7RDKEf9p04dAK7+kNvk
ci/+YhC/pfyWJFS8h9AC3vi6AF9R9PKvSRefUBemMJTaYO2qkb6Qr30INj1OotU6y8F+C2duJa5b
DiEc8DC6nyKhksnRfkkIS/nSC+SV3M4p8/zGA2/Cti3y29ikcD1ctSjb5zIrBv6+FhsVdFFbaXpl
6r/z5wDS7eri52l6pYTQ6Ne4xmdhItERXolIoJwgBfi0DTDY5rxNap5HW7oSOzwymSDzzvlG+ber
EenZ8sEmoWQjmmQXq3V4JyHNbYvpruXPS0V/lhqEJO2nGb37eyTm19WIlebrADwjDGVEb9/ysTJL
KI7tnNfEFH7a0XKMz+B9VDQrb6gBBk2Nj3L89KZKwu/AU1fCHO1YCEp7FjP1svZy4ZYOc+CKwqhj
YzXeo5ff8dG2GEmyq4hDDC/CDJT4ss05ZaQgH9gnoCWyM56qJaHgaT62JPgQ/YrG4YdXflZSP50q
lqZw64+1Eb/QwAv8GUfvbKLTLK9ZrvxXa3h9Rlly45MtHbgKXXlAfOAJf63sWiYfdR/TtZDzCVRs
EVj+PI7elG1m02iqvDw142gqKMhUM+Q3yDTaAhi/zcvZQ1qjZQ2IYL/zJg5YMFjvXK1RhVxTYMwi
gg4h59dwdrz2T4PKwSBKjOKS96CJdg8SNE6tRJv5YxfG74ierzUpBBGzzOyLYdy/bzQNJil64uQZ
1svbd0sPblUf9LdGebFEpbt94cT1EKhqPrUmgTRYXFNKjE1yJu44gflK57LKEo4phxxD+PSR+ApS
rmASXWEzOdkC7NrtenmMrRC2y3UQGZ9mrl2wOTKy7XuLA8v2DBzK4PiEDV9hohv/ZDrTahGkRGLn
Gov3yaY4zTdIzatsjioo+957c4+PEKbHSF68IKqX6jKHv82p81AzBeJgHLPBhpnGxy7PTm4OCcbb
/XpQcCynvo9yVcUAObNmaqImdRn7Rc9N3kpQ0MqztTBW40S0yoJ1DcU7v4B15AyzdBf85ONfIdWJ
8QKBGVx5WFMklfN3NlD3rorxQTAenjHNLQEq+M7zhphjS9DntyWQ283KCIVZtSh/s6NjCTJoBoXx
KBoik788QMgHZRw5zg4VOSDF7jWtTAjzoWYEyWYME9PmGDld6J+jpig46nqGGiazyGeO0rU+FLa1
+q4Ytdf4Bjcqt/qqGEZsZObIJS02xGSaWhd/0HeLawwycjAl+FJC+eYGhfOpjhg2cJeNT78WkGOQ
4qjfxJBHEJnTZaHT1ZzDYB9vQBlar8y7J5G9EXqjFxwXa8LQbFZruAQQTBsoN/hbImJELkQRJFb1
uF9dwBHtKxfNSYr2wwrFHCLgmR4VBfNxHIF7wm3COUrMpCt1omjhLdmiyfdLy1V/55VMmtSKBjsE
OortnQIqOwd1PHdSvsAYY6tyB9NSPIXCFl+Zxp3vCAm+bMB8PU3Ge58kpQm4NhD4c0jQZY8Q6FOs
+Hxu+oJ0/OZURKHVjxTFY4dcz9zzAlOlbEoyCW53ZpAJxYCU9ahWdStwmTydfC+FwsDZiw3yywVp
G/8wRenxHS3VoJ4A4nwacvjd//FnK2RBGnxy9Bdxi3+7rGEgaIbOIbXpwDiljgy1dRws4LN2mce7
09t3tTS68KEuC7ukpSSZdxwubLSK3DxwWMjej4s6gkPyoTkZsDNpn2q8VmaepI8JeBwKtdwt31M8
UCa1/V3fcxjtrQYWHPNJxdsx8TPA8p4L6eyP/VRqLsxZ0ep7GAQASElWdjgPkmG+ooLhq0hWDxvs
dpy9PbV3M4xybNfUOs9Sv4RqV/Ww3xjSLBTE2d/zuiWomW+9CmKXV6Ci6weAXYLLga0321W9W7Bn
beNXK4efRJ4iFR0QLNLWd98YmOCC8mgn0vnJVVskQLNmMoAKvdCtZ53+HOTjZ/IW6ZuzrKshz4jC
hmArKeLGHQVwU11FXxYq/2JGFOX278MfZy3r6hfEAlkD9KtIqpH7DGI6qI3BMA+TjQpGrj3JPMJG
gXRQM6JIqAxEVabJYO942Rxiyo2pbZ3dkyYp5S1xb9ZCUzMQxmZV12IjICsMQYT5f6sL8LQp3j+2
cjpFT5MilMwq9wZ4072kqCC6Z51kTmJTOSXZ1wM8tmKzI9kQ0rLrjC6XoVgiwrHLqajVTyYVvLpS
jQ/A8pYqhxpN+VVMkYZhr63BcGpZcqjdbw5oPTle6AAbJc2fdkXX71dAsLEn6wZwnq7FIXOQkQn4
z2ZeaEU+CxSATghTBvrFFFhsM/9CyeopU5dHjLRygpzdtRW5xOgbZ/fNUjLUUUuKaXmYFVOiFt9J
JzjAhYgFa+lDvc+AGV3TW7wORBAq0H8rsFKJmx7DN1dFeTXYfvuvBLrU7OwJcVzC/cTUOPO12HqX
mAxIN4s2yK2zQtINCs/UgO1NywSItH7T7HqPOMvacrNh7Y3LqgDNn+12paYDvNgRM7guSIWESjy+
E2cgd4FR+7FnH3Q3YWHBAM+7Ka2dr+EoAzxATp06LliyzjpBqpMRh4VI0sujqkaZ0kmGR1AFesmk
rIUzxV/om8m9YgI4vkiVpIoFqURFcnAUIrvgs4yU5BLL8FEbEIQCZ7QY30eHPT+yz3I23/nSqbh3
panqsDgm4gMAB5m/CAMLZUs7lT67+vNsh7HtA4WbakWkz9PjikJc520ebOHpurZ/4IlVsa6a7hIN
0UpBJY0E5Q+qeamAXymXVKU4S7pVvTpR8ZV1sc5DgErmLth0/u/Dx3mwjiWe8I0VeyaXMlf6pghb
81J7Na0L559Zjn4LFd07aLZ35oGR51HVbSWL46qKo3UwbcKpcvl1OC7xzW/EcoDYMMvTQDr2yZTU
KJXw6VfjshW9chOYoF19qEmqWv02ZXhbTAUZNhLrwaFzIpZHyQbjI/lcxBvqJ+9j7JhkLCjs3tJX
HlXutoNJhteusatHnqhY8s2pmC07zlQeikhXTmgLVwQFIuvwoKmzYs5J1hpP3AzPhb/3JxkqXp1f
OyTuiLq7U8WFmDhFlOu8U5RldmGnwzP9KIy9TtSWWn2akA5ItmRE36tDaEg1dUglRKrAcfNDPwDD
QNDCXDpgoUIhhwNGuDifQEwiVVtqzNBiIvUQ+y/9U+vmJKzL20St7MXqkWsFwOVBHnZbKWr1LbCo
oqN0TEvS+LiTic1LeCiPfLQQzNYf2jWI+H0cHLD9nMgZ22K9tPSMx8S+RRAWLEokvQXjP+3zkrU+
A9l6WYPVD2G+jr4jOROeI43P22WMf99GI9Jl5hDNTZ/7wHsGjVkLJZPvSihAqzzrmX7JpBO9Wj4k
bz+YFn8ZoRa9X+LFO57dzOlP32Zcqpg7fwK3X83qUTkkp3/6zF9z1i0fZLAEo9hHQxrF9MW1KlFB
VaZDuhc9z+hc18gpIDL0XSU5lGYGpYBuqM+XGDZ/bElaLO+XzPeWB8qZrwOFo69lO034hd31OPK/
KWiVmOfeTlDEz3LYjNI+qjLniXBmq4h39LxCoIxhGc/bvPxeRibYADQqQFS0aWX/FaUVZz5gYhlL
t0aeIQh7CCZLM4xQZy5ZYvP9Az+/sBQnUzK0lNxa8kqYL/xjMN4KJbGD++9ffVgOKGVMe9IMZl5z
ZijY85IN4Ja3uuIEAmHr4KwkyRLOdaYNCK2YNl11pFZBrm5/pJ/f/0sz4erbLNThDoG6jQJCUCQi
PY8Y6Edx9DcIjgqqlxbW5UNjgQwJYLuHlNllynONcSF4CrTIYvh0XeL5ayRdHeiqZzAfWuKWl2EV
Elrjepl4f63Ey7Bf0fKVP4/TJJ1JcEMLwbs3m0sXlJ8lWLmP3TUTmTroHhVsHwIc55OKLUva/5/M
O0ULKuW+4bX0fLbnUgf0r92RAJHfyA0fUW50fCp9MhiqoiQeU0PdDTHzZ6X91gp182I4HVmeZW4w
Jizdqm3O/rWdyPrVJeeSUhgexmh8bxQQfGOcgGTsseLNIOfSjZNdpfrrvETn0eglra9fFPZDlMqO
0K6+8HK3JDNn4DAzivmnan/XaDyMmxIWQXrLH9IWM27+tKg0FzFozFJ6JEjMlN+LpupcNkhEhkAX
FQjfdkeAhBnApu/Vv0JgBXz6E/Ro9l9l9dXcI6aR9Cuz/wc9CJCB7/+awYZ1BHa9JKTKNdx9YgLC
U4fWaqTGIJx1gWOHMX0yHSqKSSc48AXLd+huzDcCHIqg6fzfrsuXikr0vqqqMTYv84pz1EDs1vWj
MsnnDpyiOqNr/r9IDMVbSYdSCnCojt6h414onSN5W8sYGK0ivkRPlHdIFc3HQ5qEy3jrUG6O0Znn
zsJglxF6+lj96039EVdPRfacK2Q40zyhNN9D6l2krPOwKRF4b0+QZbx5/LAVXWKuvonHhZ7Cbg/B
BWqxAy/HZqFOhR/neqyDHIb4JRuPeWTYjXdes8DCdHhMNDuuNagIl7eQdO3LFbqKHJb6SdBXHFMF
Hl9DEeiZ9c4Z1E6oqJVShWT77Am3+j6/xCY20cEmwMlhJwsOOYklzKb+A1FBphJ7RGhOHJpl6vsv
lTWkMnCYeoDPU2Nro5bNltwN0xwLHESR3AYBbEMi+W8Z5voe0PTrK1Mmofu3jmTpWwbrhmqcRdvq
GA1Jc34JjgZ+cO6O+QADfkAvRSodNcCUJ/t9UFYlt77OvYiWLuDsnW1VNWBovD8ueFA5oqqBb0hu
MvLlNORwsSjsEiDne2js+Wysnpm27EvUT4acPS2qsJOTdSROCxf+VDkOyuuPq/fiKYGpjGzbgAJX
zec8F8FeIasg4pE8SkeVWmYkZKoZ6iAcBRBmWehfS1dC2IxV2sr3LfQUNsava8ZLPzYytCDigt9j
2RyJLWZQXgvaw++Ak8jdSgStIZbHjZTwTgDFztfp4LMgjNzFxQAruE59he4HqsagjbgaMU84rn6P
VGi5DXV9LMg+AALn735veZcWjT1ORPRWL0bTxmGSOpI9GQqnHTrKgr/zGz5Cry47upHjCm5H0gcR
ZUkBtzhlk+wePAdhB6PU3Lx73VMd3txnqiXUQ3ONuLfZo+egxenev7iD09OMMQJ4ySqFBbPODv6f
nQGVRr7pgcD/D3grKhsTe8Qw/NkM26ll+DigWcMTj8dQH66U9ZJsLRJtIi9mZd+PZvJPS3VZNa9u
Cxk3cld+i6fCDp72e93KP50WQfMu0k82xf8XlIU1p0XWBglwjVQvCdzQcMaW9A1pMou0f27W0Co7
SMcoH7mTZnsxl1SEwwKCVhLj8ZWkm68AnnH6O6FI1lKTu3J1+QOROvS1ajizWHE8WZwdj7pUbeXQ
Ml9JHCCdnxk33Zc2aG92BW8/ET8LZ5xLmCiP0GYgs//4bKgLh2G3Eiu1J0vHxleO9ulfZxhcYLbl
Ercxq9PihCyC+lDMfX/RV+Hj09Eb1j3wi/5VYb1xISHQIhODX0KTDQzvsFdgL3MYS9seDgz19KfT
XdB0Mo+4/ObkaocgZDUwCBDqEUQ+qvkJ2rSnD4NiSLOj3RziYQQCsCnAGg6qgCyff+2AQqRAo53p
x13ca1KIamtSBhuGmM5CyVpEKZ+dqMoIxQsR9D2mK6rN3MX02yPJPOXrfzvaqatm8EFEhaREcWRj
C0bp45li3a3hScvmzQvzaQUkkM34geNDkriuBxuB0Jbm0ngkYA5eG7JkT++aqFS39NQkAPMNcZqm
DFohCOMbtQeJT3br/mMzQmaf8gRN7p+FdImG7tRDlZQeTCTlWQRWyYl+gQn+jqO6LP3xEbWrGbnO
qyjef/9dHIsOqb0zhWVtS4pryeNtYWjns+0Z1ExyHMiKwXAy7B3vVGsMzCRL02nQp7A2x2FHXFvS
Ve7K2ChXzxQ8vPHLej8L1aVysOIlwolYfjisEMJzdP7afZhZqMj0VakU9VbqmSFSFH+GyeBMWWq2
gEVmkH2bHM7Yi/c+cTfxQBp1KN5UXUCrY1OuoSpd0Uevo2tm8A4UC+1815VYSj4BdEg1YwSjvejV
L/FUwvdwnF+wiLpxnLFDB2nmVKuVinTcdBm9W/6Pwuny0JizuQa/+BXvDf+8mUF1F4sPkQcnL3og
w1GAjjdrajVEj6mKdPMH/4gWAgwWnTvo412Hwho+JuvMIQG0BBPWRW03UZxQQ5CNG2pKo2kxIIjb
ruyZCxcjSLAUI4E/y/2IeN6ncDMsyNQjsWAvrSAWTN9ZkUwBgre3xKGmLsAM/JF2W5PLktyT1sZv
pTb61fSklylm/4w9MClE+vm5/NZjLYJljvhGH3sRO5c+MNnQDefkJv3mRqtTvbp/gC9Ri9sffCdD
7fw64POQLf18/UUSBjyw5NZ1kXxYsmOt2ZisfaOm2rOryO00bydytBuTTfO05Z4drN5MDBUsxzD5
7PfJ4vN85zhdqikYKhai7Zl13zjVtSjKyyvjcEqQyvL+HKLTR0zpKv27Se5Tqvvs3NabOZE5vNGV
tAxukiA67Hf3MWWDGi+IlX2NLVYFg6jQvvxHcUXtCMcaXDwvCDq5iIZdrOF+ngbifMAz2cdP3xcr
YBx09M/9JTSzxQz+JRJqtCZ+l9xS2tFgqt8Mm661kxcu8klqgwpJO1ryVXGMBeAn/YEC+CSZVVaQ
+y/x3sO8O8yPMuVWycamkWBT8zLATg0cz92I2cBufK9xZNmw80R0R+ChKC/pAQIVNA7CORtMd0O+
JrGqZvD/eJpE9JtggYji895xuLbU/E/QJadRSc5l14TO9w/xZ8bFcU1U6VectHwvlnJlWgruj7bs
cmUpmbu6K/k4lYPM8qn+XqpAfHFz2wee4GisL7mAsGos5K4L+jn9/aEBj42aBI03OKRNFGTKneeM
y5xq6Jk4xUPV8oGgsBZkz40qYy88V0ngGkaffBlKRpczY/RQec/kqZJRsJN99wlta0lr+uRL014G
HBV+54RqwGvjfJ8oVvdd3JCx7bZ2aKMbIbGKDpXlMgZGt8Y0Mfkbl/tjToESRQyuUlGXNPvbQJOP
rYALFco0HIfF5NZCTHv2ygQu0pLuYIIiWWv01ElIw+UcBcWpnDqJKPnHQ9ebI+PKQJaXitZXz/5w
l019MZQeElJZGeX8m045PrgxsK7We8LfZa+o2Zn/pQf2OGdTGCFta6k6SPzKqtX33goTq+GsbR2O
D60iwWGsL8u0/+ArEWDnEKblndNvKK4ryEf1jKE9wQEO0VJ5HBkn2YXLiLhTiaDCNBGw0EyaGiOJ
7scdLwEBYApgNMlaJ6lw4k3gdzeLBTDAZ6Zzeh29fATPWqUz2Pm0YXnT+XK+XSkPL9j4rUvvpkd3
iTQr8iXyKzdT/yv0eHMm4L8DNAGxiKImMeCnhkDvwzDdddoILZSbQCP5JQy01TWvroGuZr+phL1A
4DfbdUeMITTYg5j6gAswimipX8TjQOvQRBLDFOzV8x8zzvO8uN798c8cj7AZ4UKNag1QLJMkV1sl
/ObULAgkWnaqwNisOrbDSM5TogIqnhQpUwK0Y2FvRNVAxou81SSth2IWNav5Os04sXYOQc3y9T4g
XLCncvosuYFQrwc453oe+8kyhyj2uAh7CQtYPojdd9SZtKXO/8Fm0J/10Fd1R0Dr8yIHFghEKJs0
e40bBEE2bgZ0MeeTh3QFYF9gAeTBgUIZPPb7Zhsm/XZ5YRz02bL2xnJaUggMvB/dg0xABw+17+zj
1Kzmf/+JIfh4/uTtL5Hvr0WnLSIhHDeOnQ82D5t9gY+RQEBNcFvmpp8wnFBLMh+1DrdEpEAOweCz
MK0SViIHiXK5+W4wfTyxVeRdhZpnpiZAZVP1WGmWmWh09KT7PiiTn729NgpnlO7CQdce+39FMZAx
gE6/8K40m+JVMl4N7npk2jf4sJeMsUW8sD5bi8d6AqkQaN3jRiGhJAkJs/6yoNh6gg/gpXETdwni
j/tZlPS+ZzZNmtiA4l6lZFT8QrpeF5Wlbl7GdcuZTXkIaTOg+T68ZUJxK6uUmrOEJ0JbKybDiMEz
7HhXDkb1is6ZzITrq1Drx1FhJtiK+Sf4Uk1CdtQ7gsKql0oKaKE5YYKRaXuN4rWXyptEarVn8srj
MIZ3FCoKkZI7AlXINCtRcp5qcyRHS63wKcqWhdaYmejFO0TzOfT0poO5bh2o90xDHhD1ARJRWY/I
WZVMVbYySFyqBTFhXlXithsYHwgrk7SMRfnZNMGHRqnKKdw0w8lIs/rKFSxtYEfXkUbrBXuVBSXZ
JIPucBcC9T5m3607EHF/3MMg7L6jtBiTeIZxbDald5g62V1c/pcc3PQN1n/206ElhynASwmuWVDF
xOwFQYG7H84xGymm/IQafkhkHlBmAeGpkzaSus1QAz5llY8t0ymHlvqnhBDo9wKJECGkPdYYmv6D
04PrFOS6y4woCGRjF9k75ZGKXpabfwxOvxlxb2z2s+ECdi/9DksM7+gL0CVUXfe34PTz3Tx452h6
WcmHXUyZm8Vw7rDm04Rt6yr6tKeMDFmdxzOsojdIgFyoH1+quJBuyn3nsk7f6NDf3q/CJdzzTuP5
EyOeD2aAI8/KhwnmMixALh3w5EIPI9j99QOtTJ8U9R2eQSS9VT9MtuidtiOj27qy644rIGSgQSaM
eHuAAa9vNMObng6IlcU3J4ltULS+ACqU/XlVhIkPrrc9FN+FMb3r/R75nyoRPmyw02w+XE7IPuPq
GpePM3cMZlpECJeUA2vssjG0WEnmaUNajdA/CK+lu9/LLs0d2oCWW1Qp8aGl9ESS1/cNGIyXO0VS
bJ3XQYYW0mJ7YnhBJn4NzkKTAEvMwJ7SedumxwSt06KmbJ9qlsAdQv+aV2GrREAvB6WtWvPWE6Jk
8f2VomrRJ552U5LLMTBot+FzX7Sk5IHRHZTqRQKgLiFezT1+txuzvmDxXKE0JFVNBrtOmX45QZh2
m7zzkAEgsb/rBumCdIAl5cJt0eTZUXa/OtG2+2yB+2B+Y3Ip7ZHWh2kHm45oWLSz06/tWuc79GQL
VLIeCe+RigzO39fje2+kF+yjRdPs3GTWrFFx31F5ZK/Xc8PWwvm38Jxe4Ch815EtgiBrMu4qeJir
nSQnFI+Gto7TFZmYAJ+SXgcPaJzzB3J8euAnSrYM1TACnvhL7yIozT7I0AppQXbmw71/tEgy36fc
iy5rqBWgzNJIsRr3HpjS/3m8TwZX9DdjibNHjHv+13Hgp9p24B68xLV7yoVXfBZEbc5zj6/ODfoW
pCtAfo/x0A8/htRjzF4m0Gr5dKwSu4x4Z+q/msshPc0BaNpAkLq4B7Ynpr39W8WqwK1eGl/WCaD7
YsN97NmqJBFL02U1THhpuBCSk39r1TSIJZc4iW0Zumwl/1qZPk11+TUtshbrWq9gilmHA6H9Icjq
5qIBmmcKvMSLg+iINkflJWHlStYEmEtIHB3rV9zUDPLWDUfDec0XUuD6pHHuBYQpJ9U2if2ATQIZ
MkCKQ0ezOuU3lscmtHoS71FhTpdQKBlnk2SoYUCpKg8J/8AsMg9zPzY4Ey+FQpcdf01UdbnSEZdl
lH9OjwRMG+ieGMORnSES/v3wz+7+i3DuAOFOFi+h7hkhf0vk9qplz8mqysMYPZRuLNP3E8JXFW3q
BNbawXv8/Sr0zE0k8rOpXVVpJZGA5vEQPKn5xcv8qaaQQq3aS+rJH7DW6iuC0b07JaCadrG1niOa
z80TfcHV2IEiRXWgcMRO++t09Onxps+kwvDYtTKqW9jkkD/vCidmHHu3DUsuFxqyOenQnvSOfyWO
+wALDK8rD+Mbjl9VUlnupLehMQsSOlbDJcWsEsdWeqzRtSXO22XnP1Lph1F4aB5qxn0pEinDtRpF
9AQ+pqokgPbpvfCcegndqijAOReKSZR6w2uT3RVtkJEWPEcjsXr0Q/eug+v1w3q1Yx+63WqRzFU7
lk9EmbwzUZMLqmBG8QzVTPr7mYOoev8TWsBoAzCSA7kKIkeMaCeD/FQ4sAAKDUSU65tNeLeeHd4N
i4eGTLf/sspllABt5qwXagYNegUSoviL6TaAhpvQg62IIbr9IkD71cmLFA8CX937QSgysUWCls2Q
6fh7+3fgC7pKdPaeh/eNJGe7eq72PttdTcaecqPdpuQGEwgo6LG40tuukXdfpnRebBN9CuTGnXCj
7imtfCwdfAeKh38hBkBVspsmSadj6AhpAkcIflfuuQT+nOQfcx0/ZVbVlQ0vzn09L3F2q96uyosl
gSFVMt+YOE/6nGsN3xN1F1Mw3A2X3I/dUY9Zw4fOLKVkr091V2m1KPofQYuSnPzGayFo08lnSX03
PUFmWxn8WWXGrO8A6E89YFPhzSEr5u0FEDhCs01OCY/1yYd8SFZRVkXsUfMSRDiVILHjS6ay1TA+
5ketDAiYvFkd74GOsHe53hlakDHsJgzDy8ZhmD5CNwfO547qS+pL5U5N5qvDUqF5Q5LsrXlJmbEy
C0EK1mf6PnIGxwEiIDtaRW7v0ki7ljQgRtMwMcTlLpBlnC9URWLKXcvhTyqtCx2OAZ9LCgOlCKD3
yeH6kHMwYIvA/SeoABi5bfERnFM/4YrtroAQPYSz/F74ttS+Lyh0E+JY0mHN2Ms8Ngk61wd0Gwes
wrQKyo/fNjINPwqMEy907X9AkyQqbgrFTDlUzaFiAkD3OgIGrLg3FQ4vJG6+3OPBQ3ar+zGMGgjg
BK63y7wLHBBD+GXBkdFv8PpM4gxngxX8zGN4hwIGdBWwBkrdRAK2xIkwF6zabmelJFtCZ6eiIpMw
Ryd6xbscIfB8gmeBnOSWr8dUfA7kliD0w26w0rN0vKOVdB70VVUA7DPwsg2rXwRWfbLj9Kx1BF3F
e4mcKGTl1K0emL3HCD7+n7a7vOJyaLC8tKW/4HIgbkzqFnuTHBQJV27BrZW89zgIPp8ZwSl+1C9j
LMjejTAiX0QR1/QmrRvE8TwTvBwxauCw+8NddIV1hFbkGjgsB+5SkXBQEr22HwGYX7N1yYgptqGD
JXFt1YWKzJTVcj7czcYCRQ0DMHei1QfKpkxu9ySXnwBZhXM5DLKWS3rW+iTbdiidpNTzEY1EL0Ej
8rgAnu0bQZyyVhWMWG9JtdVajssDw3h32KSq30e+idUHctGaR08ev0MJG/Ytd7Qw91hxVBR4AXFZ
OL7UhZQ1X2r6SpNjI+DbZAgF+fuEK5v3NTv+LSbh34SqxIZxZxibvmTWPOwkCrHBZ45WFq+X2FPQ
nLmeUeJ7e7VL3oIbPu8FPL4HWx0qMApMpwLDh7Glu52/KegJQvnMaJ3z8W1enZpXIzIiW5HquusF
6BrvsuxqATYQ7cPkJn6ML88sr3tjIoXBZySys2sWaAPYMFHwSmRXi8WETao6vO+3sK31OHLo4mhm
Otb3K9lcKBRpqjKhZaHebL3+9p8r8A98YSts4ZZWhSaWnFrrrXU/6IO7xvM3zguNDoJsChRwa7Pq
uLNLz4BXspfA9Ea2YDJCFjT4Ph/qB9QL7ZPU/WTtwcr8yzjmyXJk+ZpZVUI+asa9FfKQoWKAfpCf
mivjBJUv92L13Q4H6dWD8e/gVCdwkDptUu3rpBzivNPX5b7dRv95Jz6W3i32rsIvf6W2z35jP62v
8Ronbn66Qza8dPpUZONCOi9xSunlZ7LaOZ3ljtAtSotcixHUIwUAf09Wb3n+o+L17uKxhnaHJ15/
elWczd+Q78ULYESYaPoZz9laC7LSTxUe6BhdtJQ2hS+v/cxvBkrDZzHfXYBM1qJXSIBxKJTb18iQ
iHA5Lys6AERmKttrWW9Jl4euzrT35D+7qKohKARSbjT091+h+FdLu60DIvFLgDG5bZpIZJbZ9FpV
xqGNn45iNeOAK5ajc454U7BpuZ+GwX6cEsBLIamSEzguvrlASh/nRt+G0UFK7Pye8sKS7o3Pw1rm
5CfSgctkD1MG7BU7seMojKdRP4YYEfSAGa7WoY3gj9vTZH8e79zk9ZoYT1HpuRZk1Z/HNkkZMqow
/8pyP0Zhgkns/q6ZakmgHkvfNtymVorlEqgFv88QaE4ssZUqozUHetXUd2DAx5bnrZlf7KjUworC
hlcMyW1PJTe5QuzdOv2jp/pMUImWdJj0uC5jMMaX0dFiVpi+5Sal/cDhz5Z5ETjbXMIOcVXojZye
JgMVqe72MZnSX6TFkntGMxOj9nNnuiIFed1KH4JU3Ur6x4LjonIXlN689OasllXRoUJNGo/1/pk/
mTfLyreQfsgyZUV1H0ia90mar15aDSSRnSJASenJH1iFB/4hzrJXWBu5iqd3wl0GPQ0f7vukb5BK
JSrPfiFwV7tAM82tX7pYeBIcWrTtdz9SG6v+RDv2ScuEhF+ZrUDpMHpg3OECJBoWXOnQM/3k2uUh
nN8W27rCz/i8ymklrRFHN9HNziziWvNMY6XKuR9vZgaP1kA4k2vVZ7PjuCf+LTNQpCQncaePYnkr
fUxhsL7gFYy9Bqjei/htxaulZf1EeAKeJgnptiVsEKRuS323ISXpZqy/kv+8208/x7M86/YXXcvS
bu+G4nxBnFWEHCVwcIOlpLaI3F+RSxszfAY1JaQ+oJgA7WRhBrP4TqRObgrSjzgB1emACbE2G7He
nyzCEwFz8ufthP9pbvmtxA45PdN6zgFI8PLoeeweQj0kjJotZ4+kSbWGiL2A0i97UjiHk/NYroSE
ZsA5h4l63Qky6U/WhCC89LJnd6tigEva3/4GiPSIC5XSS0s31Kub4FWNXcrZKraGyUXFU1xqlwiG
sKIdswoM5pNDifq5oz5yzcD9PjrmEbcIHNI4FT6yrLiBvKcKzfVktUTyXmYC3GXI49RUAnUdGIhJ
A9fSjqAi9nX8xyNRsRufLGR1nKzs9NeatJFJx59gBxUcnsXXNwsR9qZNVScfuTCaFNCLzMZvy+fi
CBjOdL2JU8snKxrPY6Q9D3PEoz08sVw6t1QAiw8Z58wIZaKt46cP0Q1+Cas0C3MnxOdcHp6yJvIr
YALNuVOkEI7FmIuhg8bzywTSG0IROR1ULuSWlK5Bc4gGiH1pU1OhRdlIYmqY41zzSVcUByKrQ01G
RLBsh+uFAhTmYT6KohvbDI41GOKlciXmIXvYylJOEZnM4GhTLWKGQdA2t1WHUaKiEvUJmLBh4VZr
VnySCYnCskxy42QwEqJZe7p9JCB/g5EaLmxk1VUSwIL/V9PhriTeFqdkmdauza7uZPv2MDD1j70T
GOrXebHC3vOtNtlMfJj9NC06GURzdngqox5wrqzdXJ4MN/zsEJB9uVWhslj7iBhU9vEQdv1lbHhs
LkPU4zM5Y4Uc4Z9JX1/UeXLxzxGcLt10/1HGEVaMXZWH05lQ7qsonBbzOMpe1QvC12wPUv7v3hbr
1ul3u3dN6YhslfQZZpLunlO8ukJNTsxxeiXhexonQjn6d6zQUZB0RW75XPkwnyDfO9T8RbyyD8W+
07nbzrwOuvWltMHTMh7GWaNddnnirGlM8KPxYjOEAsv0PJ6BLx+G3Iz4qE9hpyJ+zu4qeyTrE9nS
CkNSU91MfMNlw5+jVxvkMkIUplHmyAOGixLOxA8XPtl3uGUyVsDVX36lCpjJT0Y00Y/Cios/6TcT
fOFBfye1b74DXF2z8YkCV2+SX+pP3O8gV7xFZY83WlI92egmB0hKxP39YJUv+DMF4YGttwMnkQcU
l6MIi7CZHwVyZwiBePeIZn5V79boazDGJbVuwXYOP/swigoRrGcZur1uoR+HMpU/BRctx4BOJamV
hf67ldHf9IgUST5VPKQcy1NN4E6YkkYOFxEmywl4HqJTJ40hhdHNKVKbNZ5D4ZEq9gvdGykr2C4s
ik4KLqKTC4zmMj5px5hoMJdVfmdN2lJ0PRZCwhrZl3Caoo0PV0/Y9ZUgalOv0jf3wxeKfbG4SI+d
W/h/owoRuS2DzObHF4E7LaAdKgcthkfS+8DaFl77Kx7tQRQRtcAcZRGrzNzkKHxlQQ9d6tqGDkry
yFSYujmRipXDEkjc/4H6D/azSDQ1Zz71iycDXppc2XCvGomV74/NWsgXA4es7d+a0bM90H8Vebub
V35YeYoBuDJOTD1D8en04AxJFXO3qTaoluY44xUZ2ywIg1pudZjdKc3SbBeRrlpAFV5hc3HfLryI
FgsGhLU6D+PDL09s6GluO4s/FOL3VJ2TKZT8ajDA0IOO2TNB8AMNWEr+qb9TFHBvYl7hkp/xBEcn
WG5PzdUbHwDPaTq926BTRdy2Zc2ph9v6d5a2LDs0Pa/1897VMsdygnZgv4DQ0U7uzIvFg2Z2GyMn
arnkfIlnb2+KdTtTuQSKnh0j7zSU7DbP3mLY0SugKqBhisEFtBylE2XRCI3dQvD/YB4YX7jOyBla
4DP2zxCh0+vimvPr9s35YVouK5c9I+3qC7+DTnKxPgElfihujaIDmFK0Kd6MFm9Maogi35KXZHoG
fqL/YYuKccdP5+UG71h2BtRm96G/ax2p9I5NIWNCFjVOjwMY113nwCnq0C6//WPQHDSqS1d3ht1C
8WXkqG9nt3EPs1zLVZhPCuspcBrjQrStLc/sS8G4m/NClfdaDROMWPops5LuHkfRBLFpzpFaFpkF
rlnjnIYgebzNAvrzGwNvDrkbqfMkXG0CgsnxZ/L8i8SNLZVQlT5V6TxXdaH6kQwVQPpxwKeL+cP4
joUwF4re1OrguZuVkqxGQXzZLvtcVxB093+QBgOQnBq2UdP4GleXS7s9pZxtVnvUimQVF3bT0MeG
GWEBBvTYPeSTy2HAUmmHCypkO2WVVkxhz1PPw/hlEd6r5YLXsKliuNZFp9oZbyG32Y4Os3u+JCPf
TzMLbSWEZ6Mzp0U/uf/cDun2EHi2mU0xFdupZtz/mtkeebyiUZWlvJdMfXFaRx2OC52cyqhcF/04
ZEUZ/th4YjCc+SlWC/IlWvaDvPgOlqOrCwjZBF2HKxDttERq8ab2kLaYHBYshUNSoAUy9rLLAvkk
DMjbLLMZPxQv/Zk2mq4zr5CeoVhsYXJtloaEPn81FVqSPORnAyBI/bCleBWvsL8YlKWMxOuaolsM
FMHd53OSeUkYgdJMiv6icbdb1MVfm1qR5SbECteEbRzpUDGa9neopgKN7BdYu5rZNYQSIOQ//dkB
vbtLuRzFPDOI0iTwjm5YsMo186rjc0GtsrCbkmBI79WFtyPH6q02HmZ///zJMZOLm5bBWh39Xuwh
mFm+hVA5L+uHEwcqwuP9NDWiotdjz1/ygb7mu7gYzUWj7tfjUyeGfX5MFU+GNqml6dVjKHRhccL2
GsL6Su3XneHjEwo7ViM7CV45rWfJysQhEnUruGG2g6V66Gfoqt4YnSN94zo01WGOdMH02veUui0l
Yle85kM5EZCuVgaG9HNeBTvFtmDNQs701EUtvmp7NDds2HNvwd92hcvLgqCF1r0kHBsS2Wv+XC26
jD1hpTHLgMQ6XG2mcMabKKuXdmGQheNxRLUJGDTFQ+ZCTsBUtrap8TYMAiw2TXzjaVY30oWO6muP
rW/63dXyI4nlVjAPxJNU4BPU+3yRUW6zK+GAzQco266guBulJ17awzwp3K1hB35irP7ob9Mjn4hj
47Opdj02w0rmh5MzOIc3zreUdxGHFdan4Qz4YOykYoPuJG3d64M01yXMQUOwYEmSqlgddsXOaaXJ
kVPZbnNQS38FHPtnHDeFHWZtxE1vd0Z24Uxx8qVQ5qCB7vLFc+aaPa005YU0SoOkmhn4Ku047Xod
gLvXYuTJbXFdYmyPnwtU8/lEs8s1Aa/+nlYzSj9e8YALRsnld86a3nBLXKyptPC0RLCkZjAfZrRs
7um6mV0LjetvPyW2IHWjAc93Nn70G5BnjoxT6CcFUoTW1YuyXOrBm9T9m2p0Ef7U0oH5/yz5Dboy
aGOlw7JFbEnT0ti5RtcMeE1De4PQbE3oM+uMapYDH0hNQidqXlYV7Gq3TZnS2pL0C1gfFMkEPswJ
FdoFpPNSNJe0LH/mdyooj75M6m+nosKMWQTowo5x4/OF8GcG3ynTMFzdbczlrxOMcI4vnhy+Bb0T
3KCODklfu/u1HZqaaypJtiTrf8f5DTfixqyxTm0AKkWRSvHmctdcGEVNKgjeLeQMDCoZ92BTWM0x
ZVcKMdyKucqboytjOxh0oMwR5GP4XlgjIoUDO7epeQQ2VFJSX8bgccdjVnQJF81Pk8kINczQ2S21
0Ezj6k7wh4QYHQ29XvyasM4dE/5dPIKPizt5kWtL0pfKRrdX6bTUy0/ZPpgB70lVB1FDW0ZWeFTj
H1tinTLmIVbf0Ch4JhZ1CJmM1vsdK/s8IJyjxYhMJqvwrfYXntWSjcdVdSaDDKUQhidAPnvUnoia
gfuZvqeg8w2S1/PjQCYs7ed9D1eZ+hHz8n+Bx/YPD/PlnN5xjKPVOvac9ryfOHG44n5HWaon5rc7
Wj+xg3/DS/5QeXYA0KIppUZBJLe2ZrZqfNT9x7xF/Xw+GT0pDBbvyYHsHMv3Dt3+RJ/GhmPTJjDN
qXKd09r0nVP6gEwfK1j9xHhOJIjXQcaC6Hyv2Lq7B0zpgivNlYnypRUfOnGfsuSt8wWKe+bYdIum
62UwtH077QflrdVfErvH5DeBOB0I6CLblnOedZHC7WU+mNTyH7rMFMeRiUdxCBkMRJhTMqEuAQ6b
ZSt6QbosO+ywFaM8vYTAwENSoCE49T0RLYVO/DoNOoP4U5EbWYUDG9hQef8Di38Zj5meKPOa+cz8
VVs7HmFpZyZu17YidN/YO53Rx5CEluY+5x9HNOZQzGzNlpH+k9qTsxSUUSKD8Cf9tc5iSKd/duA+
gyu2Sa96euOysN8zQwpaJMsNqsm0LsEygDqWSeP04aERLmLDn81chzH0PrQgRFVB+9loBwSUCc4Y
GXYmTc57gYjdpYrSgTTaLVa0tdh8lpCbilqu10PG56YdarE/dsuph8pnOa+pGiL78Bor7OP40AAQ
8xlbEAWzWZiw90Sjx7+8x3qoGj3HQYjolLWAF6qjMwD/ko2nUNiZy9Q5CEjLMJ/VixmQ/NQKsJsu
/X4oRSXaXLoBW09WEOcF4n70zSk/m3Qn+NW71DYUkrF6QAZb/gI9NMNcZuXIKcaIBCz45JChQNRI
1FVZyJeHiX1oWkCQ+MCiq+UfsBz9sUt4eVniSl50hLhNWp9N+meli1RuCHxeoiifXZtH+OxmcvrD
ltu5U4wOSEqXOcxQDWBWsNKylu4ZqlB0jtrCbL844LbvSIJjbheV/KZT4jP126D4euu8oMFYQgFd
QUnQBiQXwExobhl3J8NAQeF3bD34ZQYJ+uVktf60Pu0O8PuqRFXEtpNVufBsLwUwXFLtMfsqNgFc
biwd1WlyDaqIgnQJ76yBX2qYXUrCr+nss6KpyJQsRlksJBs+8At2hCcFaQfquCepJBETGJpkquGJ
tgLVY0w+ZkFdkugZS8nkJwauVAq8wws+6uBVrKvf0TUpr3ZrIMAMkvB9w5q6AmbT+/AfZ0OskQXk
V/d3rfvN1gF3ySGxFSTtWAvzFXnumgz70QKBBYmMQdVtpFOdI85h/T/z2QZatNKAKBzOhwSLVR1G
WAxoXdZqQdGSZF+P9G5hxe26ydKoxAhG3WQ7nWO/B4IFCkNMiHiOdWmUdRR2/YsJBp5RQwJ5F86R
CrfjU22NJ2jsG5onRCejGNBW4mrp392JmdnweiDNZUSNfezlGLcG+2OfCfHJelz+naVIkiRCgp9I
BrMOPM43rnRovAjG04sXsvESGT1izxLbInhTbEQZ28tSJkSEbRMwnNVsnDLq3eNr7EMyecxAJnRF
85BxzvBWqaWMGIJ89H+AIlw4nEkWCPiavrhdLJjlZDtQYRC+80LbFvk+GwOyUGqo7RxM7jKswLw4
cxMNSka2RTu0LetoqQp+809l427zFJBppb4TLpe0w4KE/HKs5fPxj9V8yHR+EoG3G9+DE9YI60OL
Hym/sXdZFPlRrdxr2VpOhDd2ausHkSOFLkutEX4i+CAcI98XA3LS2SOIJ797P8U0W3LTzDCBNWDP
amFbwuo9LQJzsNeNaJi1UI2QFMn1g4PsIZAEKV/hISiNZyH9Nmz/Hr3YzMIlH24dRuy50gjfebi/
H7xHqaADIgf3RSmNPIUpMm9KFHnWbnsG9K0kpDpuyoH4rnCTr3JzWL+I/r7t3NxJF07DmzUDCOOd
NkO4wFmc3ymuRhboPpZS2zjH5AOeOThykMiJUM4AguYtBKKgs+sbOyHX8SOSrGwImZahajFFDHmu
7bg9LPkjDipB3BDaluK14rebD2fR1XhXsfqO/P8k8/LRttbdWWHozahivzywWCof2LJ/WaMS5DE4
Ne9gK9E5ug5loVJ77qR4kTqbfWuTfdaYHsHHYuxkyH08oYfTr6CbiY7mPZY9Z89LKsafAsuSVjU8
MlYy7Pe6cTaQFI9xhgP0Y8AOvdsF1dA03XzwPGU0lW2xaz5DaHI6/h449ZEUSWarAJiixjYCp1j2
+n2MfZ9409QM4GMTD/CfVDPOfhHGV1vyRoGM55n9R462GdYVytySSSL1ziLvD5VFMxdeKi5eboYU
1wvniEIemMlouPBX0+NEK+id/0ELB9lZMyLUNGL/OQy9nrmyIAa7RICxxW2RCe5zThTNMCnmyeM+
NJBOnyx7F5GGDbjbumF0Zv+9aHPzT6R+LU+xW2JAwEyEQZ7+mGehURW88iocI2+5nFx1TH2Tg05w
SG4X59Bz2VPOcoZLeQK/+Ri9g8qChUFEkOcSqGBauc+dEfOru6wV23JnQpm1fFPx0DwIWv45QwSl
b2XrZQOqPNNRU6x1PBUO7wQH0hENQ8VDVHkiW0nG5UoQt8+34ZTX+C23vt65EqK+w3Vxzx+2OBRK
DV5B0j/7bY1KVG9UcRbcnzMjTxyW/cbj5QpLGCcWytA0oF3Vp5/369Sy+DoC8/YTlHdrO74+V6fD
k1T/0Sir7R8YQfPx1wR6SnuItUNuXr3O5TtknPQdrvBiY/pNO+fjZnDCjuyvpCn8q3/+DM2R0hKz
jT/8fF6gFJ3di7RKtLmvYjqs31p4f/B7conhuNhy7ncAmk+tqw6qkM97AdEidxV3EDVKPmDEPj2h
neWaehV8TQ81JDe7vi7V+wEGgjq32Kl2t+kLpxfT75dQ2xNsA82Fue6X+eSpyK/6noOituD2Bail
NgQ00jEpgXMyWf8CLpmvFb80af2+otBopEXoUGH236zvKpySYabuBCYVz3wA1I3o7/fwDHQG4enN
rP74NuAgXGeqDZUTh1Ilu/GSyBj9Z7sumdamzDRvbW4gmZtgpCeoLzKaGwxklgWtz2UtM6RqUg7g
68nxXz9Hc9RuZBN756EyErebfusr2LbJreCdygSXy2YC6iB4ThZx1oF9I3XCWZ4sh3q2SPjycIst
16eD5iuDBmv2WuQi9Do9e7NgWnt6m7aLOZVi/2NHlbJG3dbn0N5iXW88Lb64GEXGRP0cNb1lQ7cX
bKU/eyrGGyyC1Ud8FZuf26fnklG0L0jHlClvzosf9THySyAFRYd2+wnfyvah/GcWyOdJggf5eRSn
T+rvLTEzlBBwReGAVA5slHafCjoKp28ZZaBUaXqErW6Az4JOV0YBnCADFw3oa9Xq92KrgoUwoxJM
CIf1wp9JDA/7+kv4YfPCwYRqfSNkqyIlOrkiSIPTnE8UveDWklevxirc8wAFnNBIigUsdx0o3ZSg
fY3vH97+Vs6ysfp07kEQ6G8oa0UJg95bqZaG5Xhh+h+OTdTRuMH0e2e4Xd5U04GdSv//qD21pC4Q
kXNtRvufnp9Atl3batPAJj5+roRpCpY/fGs3otl6lNCEVn1G6o4Em1YwzPulUU81lFMArbkSmm0n
4Y8Y/+BBUrb9q9wUxqcwgiHd7ewrU93EiwAIUJCJ+w/r3Z1RrPPmMSz8PEG9vn/VbSmcalP2S2AN
PYtdKp87UY4Vlde/dsbJ7Z5ImC8l8n1xi1VrKoReOAWaqm6fFxEdR+L7H+/xQMn9Mr02Lb/f9cld
ooHGQpPKcvVgVCoKANubynXm+0HinKI5uWhpJ/g2zweOZfr4ME3n/SzAO1SYZlePIVS820HPEra1
NHDs9jTyf7PiDYlygqct2qDcIwjCkhBRd/+2znTEFGVb3VjsLSuOczGtMMcP7CT5n1Y/cg+ZIwjZ
3o4wc0rfwfp5DPyYqeORo/0MLlFIOT94Ztk1EtkkTN9kvBQ3By/0N9IuQaYmal9lebkfaAfQ+TKo
J2QARAVZLRZaYL7hxxLACKO0Y+4LlAl1G8kMG4CaHOlsyOzsyxJxrIIPPz/YL8GDih69yhsaeX+I
0FbFBsJNMnWY91pJgY/w9pE7RrbSyP20vNtYAfpr6C8SQ+kYKnviRoa2L+2mDQd1YG8677XXaoKK
ZgMvYZHT3rl42lz/QGyD41LsQaCFW8PvmQO8Wtq3c1lN+RUmSpSBwOvyf8xpJE5uEVI7RW5EG5/l
wf9aLCEhMXeS999+O1AKp/F7uFQdMvYh7BUDy913Jsh2cYXwft4SxQCw2NgWsBkGhGTa14gh3PSR
W1i+zkNHU9mKY4RUsZrYpvHhQCeZZs3zJ95WEJzXmj5ae7VJjCneIeFztKW/+lCRs/Mt05D9aPRO
W6YxJQC9ihb4PeoL7izj55BmuzKfqhpFpabf9C520YfQ7KYAMjq6ULJ6UQ4Je3vK7LjL+TMf8xSR
8GVswbYkf4c9pgWvsvA/k0gsGqT6+OtZ8kjv8N4BsIrF310Zy76v4CyDxucZ9ZRhfdt781lsPU3u
AaFqkSzTDQpgDwtghh1rVAJB5xhG4cNXJG4Yb2yrhqY5EVWnv6rUDafYccSC/G4AJDjP5d8en/Ay
jbgyv/COwHU16ltS7sWG/XusBYYZtks5h31c657KWEwc1J+0QF5+ZmPUM0XMoya4VXaDVw1+mCd3
+7JiHV0tpU5XuvMnfRR8uBxav+2qHU/tfgSHBP/J4b+BMnFipveiEF7LT2J8wQPQyRH2pOWzj9Gf
LeFj9Dr7KS4Ge/EKyPim523VT+eZQhWn6qfWjBnb/Y2x/TzEHMBQFPQO2mEAP427kvKSD2cbZaVQ
O1x3K36VDHIwxviwTLu9iv+elGUll4r3TvLwPw2IR+kFmFstRsc+qvCG0pP77DK6E4A5jfKmLpnj
TNjTYSkm1Ti10oMCbLZHjlemHEY39C9JDuxZJewCPx9oamDXS2VOp97S2apLWu1c+lfNVTPswAVQ
HnuzjoGdSXEGDGh+T6Semp967kF6nVO2NGEr3s6LIza/p767F3l+qxR4xhCRefiCuH0o3l+G0Hpg
8n2yiE3YumHqp/6g8JBF0GrjeuTxwkJfcNApucNiavzj4WO+14BBIQJ25OrGi5lpKxZHITPe7JIK
Hfz7ga+HUmCGcTi9JUoH7HlsiT/TQG5OMhYEmkdF1eeC8IO0AaxZ/ZkJkti+QpMS07gHcJyG5nqd
QMcUxdVe5Oi6EDx8UGfa2LasRQG1rG6/3HgepJsCmyo/SVdnIlyrt7A9KDFz1rTUCdG0bjBA+W3J
9wo27VAeExQV7paPHtC4kQeekaJI4JeyrMjHuMLbRp8g6L18K98yhA/SwiOpdac25qPb5SnxehM7
j7Etm5kXqedvzMTULcO63cPf0FQpRW/oTJVFYTmWTpR4cYFquLsFkxmO8IvMgSCSgwgTMM32n70S
f6nsME8LTRpLr31B/WsOiV3jr2BIx/cS74ON24F5FDNaGQZpmXhjsHu0p0VgnZw/dOQ2PMN7YWeD
VQNW5RbSHhP3WwXr+VqnS35LeNLwYPf9Dh2Ee2OxHZ2tIEn4btSCG3lQy/lg/8Dog2Sqipil7Zda
I5FCTMhrZsESyuQcNEfde937fhK+IktgOcisObFJWbgapgPr0sR01303ca0QJOtQEPMFRh5uHrqS
gBJEcqunlHZIi66+dMBri7ncRRh/mDASUM5Wcr3+MyoFVxVCitJ0YgybQibLZEZbqe135e7gTpaP
FzfO3PgrT9/dY9dwWldzW8d1Ev4ghybsxhoxXO+8Hl4aPYTbtwx/GVCCdFC5t25cqmAWNAMgN1H3
PaLbuxrHZxaHNCTNhHU3NCom/TBEP6OnezQpyh9vOKY3o5KbbWrSyHq77MlobZtzPSCxR3KdBYNj
Ek0jigO2IFRTowQdASw9i8vGzSGnvnZaJUOa4gCpSfAsz6iOGZIufHGXhXABgkl2g/HRwyes/F2T
x9oMocx/lCyclUUXENaDEWUGWXXN7b/f6eJLdXXPMK00LZvMZQ86FjPXqiRawCDn5eZ2bKwdwiLZ
KOcrIREXjCQbuaR61Bvg21Fc6O1sycilHiyIdIRGvgTuuVE7eQRyz0WSNiCN0TE1l3ioPneT4rMN
tA+mQB/Zbldt8qY8jsECCUAOODxXGqQ3kkKtgCbr1HjMWqbtIPn0iYm0jwY1QcJbkHkkaS2MK22x
jWvVXS12w6nboQwOKR4+rCLtwuZ59CUrUua4O7Se4R86a0hFe1rYe3jWMhrk6oF//lGwswMg86oD
6CWpUQpTFKKkxm7JGXucFosZVMauc01DrAZOQsmSYzpTVIet9r+fDY4vS5U3fW7ybDZ69L/SPn6H
p/DOsyqFB2KgIZxxUCutR9yHaFpTHZKLDWXRMXQadn2yoOMkyZ13rd1UnA52xn9WpoMCthKfkNMH
9MpYUOVEElrVEbzP2+nNTn3m5liRLLE3PIhZdqMmIn8oW8S6WQ1U1mBSic/rU3rxiI8EkG3Zm9UM
QFORDCe2XOts+XS2uipuIlGWpi9EfwEPRSeRLx9nmY4lgO3fTq5D7i22WTtTeW41thg+DMJvJdnW
J1sKiBvo3ku5c/Q/2J5kQ72LUsQuCHtqjzwGIX7rhLCr9MT3tSBoLfuu3U535FXpdJl2c69+sBDt
mEls8VgT2hf1x84XF/sfHtOU7JaHqda83Cz15CagRmsg1RF//r6Hi4E8J+K9eIUxm7uNc4zdcMp7
epO8JYCtKPW73ovwtxOrYVE+ICxbbGf3L/ZFRgUYZBD9dK0yBwsYvRL3k7anM6MRDIO1HqseWh6G
OZV4/lU0mmOmHwOyr7ln8hKPDV9wIuN7o15ETuP8FoXMK08HGNC3WKptCoeTKLXMko+1KRuYRX2y
5BsUfTx38aEXgwsldjc9dP1rAkMEkHNyPD28i5rjwATxiwE5qWLVAqHFfp546ilABLEmGb9OyA/Q
5E5+nhSq+AtvoAnD+hwMffAEI07Ie4P5CaUG3D/38JKr03CFU/7mGXw/U4OleYigLEwarzUAjwN9
HiwC4bMl9wFR3NVQ+kV2pSLZf79xqoYjDjp/zeLPMupZEgytOeuhIvA9jbY67gU80yy63Q5vBZQF
9EzvFJ8sk7/BVrtVlgw8UcwvyxG5tN9Qd8GeT45BHFrvGU2hcMwWVihKpo37cmgCztah7R0sjxKS
coCOtiCuJmhAtZuqOJ/V33+N4UQ4oZSWxGRYcD0WZxjyHQV0g47gVRi6AUzzY8s0TCnOQs3Md9ZB
A/WojUrm/xorAVTRYtmNJlUdz4mYDj8GOJro/DF0SVuPcHyq0R8pc7G3vCX6GDve2xAQWFl5c4++
wQYqNbwhssZvDAus0fsKtHIdd6X/op7zCbgoV2PxXGW5K9nBJUGmAJb0XPaJHAxB8T85AnD1yR98
n5/IXX/qhL6Z42LTSPIVMHYnND1F3o3ftJ0ecIK6jmV9d8H7E1p1YB1VNiQrUQjew3JkBOEkbQUM
/vsVraAExk61cRXLfpUoTvJlcNY7f/OcTCP+sTA4r2Y5w8UUEyHh1mDcG3itSpPKjf94h7NhBNgn
Vdz3RfhXkaldLEfrSa/SKnVE8lA1yoxme82HweJdnC/I9CQtGBqADx8NuSkPFn+570T8xz3JjLut
Q5wS8gv9JWHYTjI+IEFakfG0GiVu/e4WQHXhtlhCVMyKZs/Co6VARDHhwBC8UGvI4yC45d3brWUq
lhzcgJk0/3Q4UrDYzvZqtoPPMmhasvj03TmpfClZzL7g3CUHPy5L8w+0OuAFkhdX5IZ1ZN2Cu6QQ
Ctg2WxaluZO30IH0BWT6tIwhmJn4VzIig3u8LpT1ldaecoEMsQ2jxOi4ufWAE/smuvxdD7/ZVhw/
swHxx+QMrxey0hfmL9vYsC8O2Hj7z4GUTvuG1YdGszP2ANRJWro5X9gWC5h9eH1WTM7rXsQqFdqs
PtI+RGuZW5q+E9ymibqmt9OVxhV7LzWIp4zySXhzWxUnrZvEkcSL3Qqppx8NfwW3TFpfLHZARXwM
vQtjLhOOYYQ5bSKVal1D+gfyiRjPB7cCYlWpZo4j/4f8cxr1hfOAIVMG4iVqw0N851MkTufbSmST
YJUXF/yF0aZPhzKJxUK+Qmn7/Nlu3iiuChVBQiAHY6jGDvEL3lmZtzyRLkVK80DzdSAWfwQiL8SD
QNGS1XiBeDZDCGgiyVP0LfCMvn8rrAnpQapYfUo8cVofBl2S8pIsSx8IoKBns201tqFXaF4Zxrr9
CJeFFrnkWUSTvFsvMHxeu0nnDlvGyvinqRaH846VLN9FLcYIah994Fvx4q3Z0Ba/nOVrHk9nWHfj
plUb1a2hF29tleO0uV+uprrx6jwuyYKpi7DfYytp4SlPN0AxXQfvUPcveaHFzwKrVcg3+bBAkAQs
KsBQJiXlnjOk70+sj5HglL+Y1UTNRVv1bTzIRfIinXro/muq1URTvENyaDzIZCEGO2kM4n8gOV/T
NyLADtpTPLzWD2/K2KFOKRFoaHgrMzTe442hxl7A3DKECG0qcY6oW+1J25SDKuO1pilBCtA4rwuk
0dNVmypBW0qqKtTi/LoOCvPzzn/oPXzxDHm8sI5MxEPl2S/Io/zzymlamAA7XPrSN9ct7V5Lg2QI
41L8NEQDbvHXwDXO3rHL3bvp9u6V2Uo0nS2RDr6R2fHAxQySXx0p+8VqvrW6xlyhw20mEX6+f2uv
ojcmdUMOmfJQRhokNuoZdf2+I/x+eYQFEO/n5mnIn9FZRZc/7EK94QRKo9Omoe1VfpO51JZ4ojEO
I50qE+eZSPNusJYbqm168VC5IuSr7U36tNinAq45UMKf8+rnOOj/iiA3/VR4cQrJT47hQKYrNEjG
dDQsDiqLvaQjewuw4tI+egtowai2a4Ix1+fbkyJZHBiM75JgYWK4c4ZCj3Ae8AoRSxUMo/Dcmuvz
EYlzGWJuvp1+JaBei7ON/bD8mdY1HnjuyuecJ0a90qtK81H27zf7gpN2o3U7L9WN5+Xib8yfF9yq
IevelWacYVVjwF+CRnVV7fyXnZ1wpt+C7qfZ19VqAJbILt7jwbpXfMloR2GOwLuUy6GnMeU1jyae
gKZ1EDVpo7FWZbQSjZXQVrvaKOkglaAdrz9pXmFEOfj/3b0lUUQMT97p9/Y7oXUNnekBE5qCQm1N
ys7gKuOU+eLq+vc1SLQZaRnCha38oPvEJv8/VqvrmSKBz1QH5oLJY6KH0zfh7OJk9VyNktT2C+iM
Ngk6hvcM+SZ0kdlFPKzFJ0Yxl50d3sv+0K0wWIafGRDEbet6GOWFFusXdsNjnRopa0fn7atHezo5
cVomdACVlvgfzDs3UWEfX5kW5oPXkggxgNm05K4OvekUB0qG63qpCjAgagp44WJCvCHhhS4kr3XO
zI9SWVoyldQJI2iIZ/VClXb3W5M1oSB4/GghuvhYNESAyUZEigxdh1xpxwTniuZyvMZFegv9n2C/
0CtWXuvQvXPaMrKveuEPTQ2KGbbVNKhhaiRs5qvEqFycTsbjacTUntNomcpvoq3la0WSsDFOo+m9
Ol8gdG/gWqY+9KvfgmZ6pr6W1syDvrY3g3HiSDkfvAXgaATTCdPKxIIkzmdPk3PFxhP3JcuwiowM
+F8gmLRbMi+8NUE6+ZzJr6rVdICSOcWhtIbhtc/5my554xAJHsCsLbEf2EXdilH8P2wa76CLKoEv
FpWiV6PtEitIytYgsGmXyFW3cy35Ti9qxKHPRXbj6KnU8KxE0C9ZEOZ2AQJRPRgnMq0zBtacHASI
BHQ8seY44HZEMv669/yghnDRGfoc1YBI+FwgYlkff13tVjA/sETnm+SBi5Xdeail2Esfj2ex+/bC
MUOq/YYhhdqYsaXCHX0LYuznh99P1ZcvOeHiCycSxZp9BAgE2dE7IZCDG7LoLwGu+Jwjm93V1zgR
PqpwMg+tDLiXWB7mEk1gK966PnoKqgpprEVNClGoE07ICp1A0adQivs7dtTs6e12vQSQTdepPgFH
+le0GEQbEiugEYM5j4zg4BC1noLh4pNS1TlAxSyPRBrbrOGg2rzO0XXUJql59PuwDLcqC3WafLgV
hbMBDSc7hbJ+PfKrdjQrk71yRx2l8KhgIBG0H6F19mQdJagW0VtrN43Q3Rwd12tEnbKXI3KkOPCR
HJgTRZMrEV6lfNEABEMOYlWbXbADCPTsWFQADvkDkhygORmkcCNUdkz+PlOjHkM1aKfpkQldek+1
CoCDlodfWlJrJdX355fh7ROS69Qj6/hsFmW9CG+w/8+14bf7uVwpyokpITDet0QVjDiWHMG4uOGZ
IBxfBOP4ff4kn9GmNP6nQHhyFJgj83Sh3KSdZjgK5cSSwTYmjLg2o6vQWtdb8lf5VoNS43YSgyQR
p640dsGF2DbyBopERIvn7nw9oloW/IuuTPEg83J9ar0+G41DjWiQLFbKss8gK+OVpldPCjAnbfSL
ZTy8BsxsF6NcxfBlN6QSTpM2NtLxCOG0WGASdhBEjPko/hGNyAz24liOnS8LpCa7o/NbPp4fXUf6
1KIP402s8Frxx04LD2dwmPrI3aWMeYerPaTllreo939MegH9SaLt/+ysTvPRcZq2ez4p+RpAHsjb
ztrknFky6cnfobpQccK050h5cUp3C8vVt7Z5lwJXW2Hl/cU3a2ja0WGettPPBNQq4YDY9AcH0Kx1
Qgy+O5tSiq3HrjqLo/olxGXSUchBuVVtcV9sD5QYzKKbGHMU7MUWyvB2X5Pw1NA2Mn1WDxshvvMa
sPAUekMVyD6fAV1J2e+7rJUb7EEqeBjoqHaCxvJAZWtCWB7m90ZvrBRl2IlRfcDZQ5etoTLwLk9q
fmbcvaD4kBJIIVKKbCGDa9/wQUtyBa1Qg6ynP1DV0R2HwZbCR9hMxkCBnH2ibaiv2kKXPrYqwsLb
uirja2vtbNzIOuwyHgcMgPt2Zi4GJe35HcMSpsksGcYeYs86SiBdf+LCiBzZxvB+6K5WpwDKS16d
QQ/tD3wmZ2ieT+86u44/8ukFBWTaRJZJljIw8ZVblZUzz5cAa6wbktgrO2+wnZaHz9+zXFQX4kMT
/H6GvyWdchtfoA0FEwqkW31FT2i4lTvwqW6PcKPMpfvLojx7AUFHGMMjXDtMiAEaPAI3guiFsw1+
b0SnkuJzhzL47++xzh1IzFsmDMnU1igW3ilCGI3FHwYMV1FJG7jp9l1To5NtkQveF0/YAZY90hSU
yxD7mWYX7fHih8YvD91mIFMPtGTFiEsU2R+b4YBCLAQyf6cUYRJKlY9XkHMki/PmrHrM1d9ePYWd
qHFCGvG/mbfpT/4ZBg2Sclocs8KH7txlqIUfR+EeMioqz2tWEJHIpribnl5X1RdrN9BI5d9l6Dl6
q+cyyEG85jcajND8EnzL5h7RJgt2V+gIdc4Ajv1/Dbwmv4OP0GyrBuvU95eeod6Pa/X10+DUpm3a
6eR2aSZgECQ8ER1cKmo0PHFYkJF7AGT8WeuVnZgGJLIH7x4Tp7TRbH1Vc5BqQfOcsJEupgdTbcjl
RfnmHrCu0ZNcrLUb6L/1hgWjhLbj5Muo8ZOCsAwhPTaT8fceFgJzrrMZG6YEiHmexrX/UsYljoGk
hWkw/iKm4bxNjSijobp13cAGWBEfPHNYn2rXkoS8Gxy7GInyD7RYsR26yLRZIF+vYZNUCuFWYvGD
HbRjdVpb+nMadNulOpPAzrLVTVULdmmqsQ4chA2p0DiCxviNDTD87C14O2kDjZbHXmkbZ53U/dft
vy0bouzzU+Z+OOGTHOwvqe9efBZUKuwee6lEZ9TJRdl7LAhaJOdzdKv8qdaELazb83JG3fMdvD9j
kOdjtUDDpBHPVpwgQAhTVC0qiMIUCQH8NbZzQ51fK1gs1mzGCZm6c0KpgyebegCS6+2biVa9QikJ
DvbK2iiyya5A1bu0HKs4yTv4ncUEdtgWnBNuTj5uaZRjhAODQCxqsSjJ78DnVbNI2GiHaJs8Ilw/
cT/9JjLKHoOxbRS3N2wV2GeN2hbzDtXo1q5hPeFlOYMtAtXWLv+9XpNEvS8M/5+tBjfpBYp41xcm
cZadKR9KuWPOA+nTFHWioEx4PbKjqFQ33yzsXHrhAsGBfc0twuFCfXPeHCwoDd2cmlYvkDSt4NrY
pXrK7fGHu3sweYYf6MvNiflptMzWrnEPkF7zMTtv7kbMEPMzeGRm0tP7TvI+xG90AJi/USmbv1eR
r520xAJWPIMLJXOMUw97O4Vo/gJ3bMzL7JXUl92NMLGFY2wrqVKzh0/L6rHBjpAu8c3nR3Zvix0F
dDWndnOdEIVlf+orRE1vL0k8y01UY+piq+F1ilvOAkhz06WKVbbiSLXNsXCAbu0CoOIEoWBb31mV
G0uz8Dao4H+uwjaGx2H9VX+dbN7ZI+C2l0jfnJGbBmJU9XC2U0PsNHOque6KUhApF3yjrBlTpJXd
XkpL2bKKUMGgSR+AU6f3RAQ2krvFTnLPEnaAfAeGSFze5GLoZoBzv8X/c1bobZv15fbBqL4nUVJI
Pk3vCMjqNjZY0i98BTkTcs82HxpOZOB9CUvjVIEthpbeVTZeELTIS8j/ADQygO15LL6qaQljzk/s
5ckiy1h3pj8x9V4PiAqIs4GKMI7bG5d/RT3VvTXLPeK8sBRvX7WTxuADPI1uakQqhlvdgdynmLIZ
oeB/CpGP3ffkpQVm5TverxAWStoNt0j1OB6OE0Ae+qVSemNLknQ9yZDzZvLmYUhhUAuGKW3BPnN/
PolcnRHu7ooGFm4/nb78rxRQGYrSH8Sy1IjEk6W4eBcw5HBk+6Yd4KoJodIb4kwaOrBGJyte3J+n
3X/PMMM9JlS4aByC3IzYcUKGgENHIFpihGEHo8hzLuKlF+Skvuqwwc5DpcS5LjvvXzJiuf6KHiI2
29K9K9n/iLDkn7cCNMV1Lt1xbFtFWnKdELURnfyq4ONBdPTAE9g5sikYZLihVjSSqX/pA2iCm/DK
CbZxaqcdIRCuelwjW7fleNKK6Uea0IrXxizB/Zlrp2u5HaqvBKY6Wyiw3A7x8apJof65z+MpvDzC
ATR2H6Ihp0SuWvJIrmSr+rwiRC1kX58X/BrxvoU/fNWja7nJZf7Sb8uPGjzB4D3CWi0ve6MzdNhY
gF5Ku5hsDMqddTxu27tOgmnDvn8VR6HQAZzC8si4DnEXVfl31JIHWm/etRA1KuSnPVR6bNKgs+gs
0bduutxo56+/mWIw5RzjPFuvjuo/TzaDNBOW/+ofeuNOFXNKvWHsLwucrUMyPwbKEwYqcNdolXS6
u+N9ouO9zLbdN0fPqx22N9n1UFp2jnG07UGqxZDehjzI12gV6TVzwmuR4xPzPQ3gyuzlBBTCgniE
aOdh0nbUBM1lOTivo8c97jlWaxWe94NzBTEMLvQuaISpEKuyHZ8MfjunBJJ5eLTtE8ffHKn1b3Uk
whF0gPrtuLSxi2evLddX13c5oM/KY+johz9++ABNG46sNgalEQmUHOXXKIj3malZJ7qUtbRVLk4T
khf7Xp2dB2APkZv/zk6mZndK+9pqh3Nw4tSd63/WXgShHRrNlNlvHBeFVwXVasv5/FXPO5xLwlZF
cXPhwY2zhWqPjTt7fjB1KVFxd3EFkKqdLQBDvXXinJ8+IBUGDsjzsrO5PqOItTAZODR2oZYj6UbH
CWsYTLrWC0vl8Znn5N+eJzgDRiPGjDs51kQ6UC7l6CvFrIlcMnb+XK+4ZtdszVEqC3a0WeFVv9Uw
8RtruvLYn/xVEm20C8iiwz9IyVmQ6vO33qKXlxM0F7BPkaXIEK87cq37zp/Fomj4q31lmbtENz0Y
BqouSuWhRnhZ2VjDuKd7ksPgYFzBEhliJqFhg+ibYdKkB+nQ5X47hH47v2M1eNk7XvokPnCS2xI6
RC5Hg791gI8NkTcsp/3WK+IbAjuvkiSzLiRQ3Iv7AQW9BFyG5tVFML/ZlYO1mgDYC0qUA7Dbx6yb
cHqX9m8BBEE1GkxPPt9ol4bCOED9+NME7d1Yov/GqG/n3ofYh9jMdrvtv3Rsi6DH5S1fpc5wfjmX
n9XBfBPJhdoTFsx13z9mYjrZB5zT3YV8rIWj/MT/Ft8ReKHtaSMfoZknDXNVP2duMqIauYLTuAg2
t+IyGRlqzclfXe1z4lSNlykBfT09qTImQG5ovxA0xXemCZgmS+5ajr+8H/tZiIKOhoa1msOXgY9e
ZMfc1rMCOmxBitPeC1YRUPLQHWcjMeXlO0XQqNK0wd3YyxJaN5g2IvdvFY31/hlTPxL4ZJpr271J
jz0AiTOG19AQPKpZAhKNHo1008TcdDdMbBW6u3Rsf7neQaMnodsgCBmHPAmJ7sVsr1yGvCYKDlmY
55ihKMl8UaAcpoaXQC6B/H6rKHjSIBMESUYbGxTWqpekw0mjUvd6d09QFBcT0EMHPbyk4Jcv55r2
jOlWsBkHdgvzruq44QURF1WMcD3tZcma9Kx0DIgIyrWJBZD1lAHlUiGm3XuT0AN6/3ZOOGvoeFnj
YGVjcBwqLnortkWbN/Y7h7H7XPFrZswx5xCXWUuPwtL36zGHdV0/FwgbVVN8Y9M9YCSy/MerfIPq
bGCkVNkqO2SjYIxi7evVVH//JTh5tzXZnaWWvf5DATWHtRfXjIrdi8gcJEVqPr/lYyr28Qw6vrpU
QnVnjQB/Jl7+qk8Tq+1FhVS5kZOYlZS9us69qayZb3f03wl3cmoTyC9LAIobidX759yomDssIzjE
4xBXLlU51yViPVUSQZNdPi3X23TQIG61ON27hCQ5GCPrwLBZcYGUGdPiiC4W3YlPe6LmxRaSSp66
+RE+sTGGKZg+8R8DevEtwE+7MKR4T+lxJ/mdyU1NeAEnpmxOTGqnmDIzwG5m7P0ohFHEMt/RS9lB
dKj38iTxhtjZWuN1WIyDbgNSWBAIpUi56sRGD42jCk2sr/YLOWl3K5Fc+/SdM8uFpt7ZP7PdB5ZE
fQ7ZLD7GKWhPwIc9LczWypUB93f2QYVyAdhDwOFmG0d2pErEa9zAFol16keEB7+gnZxQ2o+vDjv6
5LVFrPd3I+VFXtjqEwK3nTRawQDyZWI0eo1iMf9MP34boN726la1erOvrHW85dUdy/7ZXS0RHDMS
xHNRSP84P9iPjCFe+kD1jbcw+hOHJGKf2TpxkhOle0CEPKvueSG4ZEIK4gYvIT+ICHvu7Us1CDR5
Y5Gy/YIqhAe8v8Uh8dMKEzPasWZhVIXp/oa0/klSeUFNwzk9rfGEzDf2eNbz5DlcZe4cyJMAmQaZ
t2hXWePT3TQ7ilCwgIDrMQ0Fw+JepgvXR7LR4IfMV9VtLWBJ3LjVQZzX4DXGKLyohqBVcHsXxYvh
yEpfELuP/SESGC5mY5Wp+ik2hoRVGxgtRtIzFGYVoETcM+q2Y936cytAE2Uilwzf0qPa15Rh6Pwk
KfA8lPWOoyb/Jb7BbMjkfCMq9eP25ondyul1XBWA6aIamUVz1HTPTTP7B3j7b8gztgJ/Q+zKI2ot
ykt7jdyy619KbTP3czh/6dZ3DKPgHz6YN+Ynz9AvNCB46bP1gqvEwhd1wxGpObJZD6voat3CNMQK
xy+eFMWkhPOdGurzkGrFdI8SVzTQvSG6/+uQTUB0Ml1zirhVfQU73nVop+7qHLR1BUFoOooDSH3o
iiBvsiz9+5XhZiIW4RfGPsZh8i3RnqysxxhY6YrvMY7xP+aUNv/6l34D2bN5fy7cq7wEWM/u0p8M
MHMsacDBifPrG6daW3u9t2IY7pzJ58YWFOw50YJr7Rfwt1G6CkgxzOqzrYFBETyr1I+p3azh4FEU
isIHMNnVHNgG7EsCZssQobRvhNxu5pbE9MHcboqR90D54vSZm+pwCdktOf1VhpL1IjhVT3jScIpi
YDXT7klX31r+UpbGp6WBWQ5otnVbvJRW/xihkvCTqQOHS7aAozdM8ksqeRWh/d2YlT/NvdJ+QBtO
Hb4IGHhNJ2wGLiqKP+hrKXML4ubzA5WJphNTgYKIck8BlRXIncPqjM07IOxnhaMUDTgTqX3FpvrI
09MXi3itLPPRxQ/LAxUXyfAfolO9KvHNerksfRJIBCR+BDxd2Vea4DTx4TjcGkLAtNBuJknafOu0
D+KdAm6zpoNYJU9k9Z8HYAtfXM80kqHso1nj6H/IQA8URG46hvwmPYp07yZmsumbdyUZND67eKh6
UL63DmGhFkDJdJ+gKqfQJgse0bRQHE8F3GqfUT3Q9xX7kwIOx10U57N9sUpOmBpvmsQvDjyGfle8
b3cT+/xL4tXRZYMFuiyE9tK96uYQBAU4Yw7TdHAkT1abkT8snINilxSybfvGRJ0x7OmhrODXScQW
JErDQlAeEfuEknOrXUoL4kdwADjH4ajOL6VSVbwE0kjBaRgB6cBMc5p6lyixAGgDNkDRc1vH8x32
3h/p6kylCMs9Fjx7IgjLAjEG/ekLfrxIfIoDUb8hFGo4xDb2y2pHN0L/6PSpqXwFjg/Hq4toWdPN
q01rrwKUG3idovKxjyn1ROOa8lrL4DEZgeecFWjdQjiRRDQFBGYyGhg25218DwzR04527MxpPlA6
CRBPJz5/myp9+cHTo+D9Yyi6QHNzlS0WYuouxw+dLPbWbyxangYbZTz5je76/9ek2P6uLfwcW7DY
XQSqPOmXx4QZ1CuQX0aZAQsBG1rhd3YUQJYWJjA0kX0Gw5z6FX2QQMtDW6DInYl1eF8HGSFBJmtV
D0mSRA1EcoexmOKUSsM+PcuBo6vwePyTOlIlwt4u/dBdlTyVSr9Dq9KAblNaLtPgFgA632+3rFaz
ua+ycR1hYDTveNpzALHriGEtZlae2S5x1FMw0MyYq7NhuOuPwqLJvviYxDXv8z8hmLoCCGwW04JJ
HOSlP4ZTPOAzJsqwLS8Wfr36yLapDTU5sPblR9NrYPbu3birxNhsyayMQQ8t6nBDeHrSiALJwy8f
Jmi5A/Ry0gPJMBIUVwYTgHTEwUVRIgkQ449mUFBqRQ0+8o0k81PLZeFOtKHx2tuYG2akaD4yAjBn
rWfVpMhX7favz3O5LqQK3R+DbDCTVnx+DkG9bA+ZSD+91jO2244Zy/tipjPQnS1c0/PumKiO3+we
cAK7oCVQNhHj7fB4PNoAJbniqeFsS8fsAFp20tAKRnIQ5t7mej6U9Mzwj+4z8RVBowkJK5YwKitG
Ju1vNKESfFFlXz+nmURHfRkufiPbA4ifrFW9MXI1Y7arhlsriXcZR+4fpA8Lk13xYXer16VrVT/v
lsdPWTBSHsRCgNuReL194ZWn+vvGhG2JABFK3XCTXZSi37CCO+cuHwC/2B9M+u7wvJp5qwm3gpav
mHJ0DOFR+pz9vN/LtbAZGfg+pc4XZX54MBLXkzU+y0uGVNadt4cAYfpt4ZgX/dZe7l/AKUuTJQQM
F6ZET2uQgrYYCYy7bfhtsk61b+DDNGr+iUan6xQm0suh/0pjLZuDTAENq/edcez74fo6BE412G1c
HxMo9uJONj0ndYFxjJS7gz+D5e2S7SpAyeNDLkOLMUB13ne9+kishyApoHdkUGcLARpDwcHtoDtB
wvarjIuT4D3jxN/PdBIuN088pHTe1RpsQLW2f/VEWZYsTkx1yAuCbj5lNL2TMJltYDRxp/DnP725
XTpeTxXcdGxxTafBzsVh+VyIk8SzZVYARdhOp0434Z+KowqMb6zxLAy6QR8CncmUanqHO7SeTtQD
Dd36vtf2+fpgifkQDtCqrlGorBoyJTi92whlLluYhknpJwIhWTVMMcXEgh+huVD+YidvDRH3N/8r
QenWlyw2WfFBOWjo8BJlf6ficfhWYliH0MP39mp4OL2oSGWHINK3vmbI0gTgrvi2svvJuKqYFcEc
9atI2HR0iAQCia5TgnyUJCbRxp60iM/zQPHEWi5T7E8kgNLhIy3DaHWdDK1+0mNI1It20ox8xYRv
cae+KDro2x4mLYGMredM3JwsGHh27/Str5ApPFaBLhVSsOUdltpDKH6l84o1O/6zDoV44ddfvO5G
Jw8+Cw5OqprRoH4LYB1POzUABlFOAK3kSZu/AQ27ooxs63hLgwYXR5UqQ6e+KwUP0ZJjhsya8Ohp
+mELl2T5L2hVHBWwQJpOU3ybbGC517oFsdw3fEaGs/VHxAnA9F6e0dXsTSwN5ACrN3YRx6JfSZmZ
D9bBPRAnMd9JzDDDPKb5EB8iIJob5cDMbh55+E6gn/9MUcsN9oLqAJj/AgDL2lK73QwGinykwpcY
5d+S3Xxl4j11gVw2mdubFe8iIMgJdz28dDZsg2bok/36kwakgtX9lWY4KYK+qK9uLzokIIwl968m
46ykoJVoYhBBfURkwLhCMajr5jvyQH2LK9daViEt826YfM+nag8LUrZKi8z/mP16iw+6QTpw0nNR
+Rv207cKkcCXJ922aWYcKYCQSyRCkETJQU4jnIK+TQW1qwANXwqS2rB71dC3Xh5zTtwrohTd7u4S
alTr1dCQf5jHEMqf5Ly28BWdl9XGAGMHzhsFS30oXNTJmUVTg6vHMj2swFVPdi45iEMV4pm3c+s9
UeVIyh/obIlQ2m3azjIHTCRRlkoDq/6ANpNtmBYnfYNbHcUHBSl1v8CRsKkxY2ThoH5YrBW4xFBR
drFNyM07umqHeGH2DDcuLx8pJZWuOR9zWRl/sTwHtSsauUKK2R1XdW2ifXZpDYdqClWv5bePiX90
auD1yEhdG/IaX3kwvuEUc8EkoHzDYAj4CCWP/0bwRI/kKY76ypoGGwmfa/XIMNVzKLie79IhJBOR
HwAvu996+QFH+drKONiDJ7I+A/6PlTfAR6pmbZcXA9jHaBp7abIYwkBWmnv03HaVT9MJORdKTJxT
XaZND6VlzPL9QFdZpZGHLwyGZ/smWL227uURIIqzH/GtSOcv73xUYuA52zE0THc02PoIDqK9+e1y
wuX609T37fs0YgcFBuN/aEmyho0yOVNPcQsTfJQO2kvEJdiBD5e0D4klTx38LIRYEQoNU0lQmlWc
8cJkttmPeKVAfDlDBLLlUs9XnYDtKXuEAm9AmgiDMZzrahAJZF5+S18ySaUYcbLsDup8CBwTGmFf
Q6MVDw8awgQUsiXqhhs6lVFDwacRrGVx/V32LK8JBZqXSH47NvH1xmDVC7ij9ofJKhCUfqHWYByC
bFv2+a9VhbM+bjWNNmJDp19VVkJY+Vdul9DaE/I4UgzufnenSHm/5ZfHsW5EwFPzqokhv9DA5+2F
mstYYwDSTOMvq/5XcpZMHQQ7x+cNXnEdLkpp5jgCdCAelSZSshr4nDjSMsGDNmTxO9XeO107/5Wg
vVvqEl34hKr2T7e5YrGRd1tTcC+L4UbDxDHyBzAFzoylukRf4YSKJrrGaZfUROPqFFAuV/S/gAxN
MY+GDdotdNn1hWFoCsQunzyuo+mlRTlYmx37FsWxpTpmTnbxDzILOs81Xh+3R+rspHQD4CqpnEn5
Vfft2OyxMuUlXPgMuA/y/o5FQm9a018h9Cooft55f1ug36yGx4J9tUQPU4F/Rf0B2XevQdWpKVpx
2MfpzgmtinxASL94AhuWEyeGqdatCtgne45W5ftsGoyn6RkGCiJrxzTl2fPRyeU5sCAnM0bUqUau
NpkHdgrYM0xeQrR4Uy1FDSRGQMmx/hEGfIEMm7HLXnro+Z7VV8ikX0GY+FrYDN4zws6sg6wPv5Mc
Yw44L3qRX4lYPRNTDsS9pqUzemSaxmhHVvFD9n8pgxsXDV0XZaBkmFIYTztOQ7QW/dKBOk6WsQcv
lbL5dJRcWAncrL/N7a81PWHEwLXr19vOgXpDqSv/dz+KLCvBG2+vvsuBygmoBVo8kffKi30GcuTW
lJxWTxJi+AdNCLsxufgMQZaOHLkmw7wX/qJ3AGUQVpYqAKfpHZSPHDcyeVs22qSK/y+1H7VN0UJL
VGZAceYAjdBT81urVrQHU+z7K3MGotkT6Ue181mRdHyLEznnuNjBpf3cdwAqMNGyO0UAatHpOBYT
uln4d1AxNMXFjE1nDa67shPI9Y4O+fMfBw62ATvwx1SxMa1ZwhvSdxq9ucMRQYSMzjbkMipq7lv1
yTsGKx7X8DuEeZHhLXIWQfA9mzajmo3+giUAE+JNlvi2d0ZkDmPMOQOPVrYlQp1uprdkFLnRpiRP
zX8bVphj70u4q5+iYTLpLjUJaSo1OFCR7JZf2+KO/EWzSy4cBxON/RIIGjtPRG0JbW/+IlNyNwRw
AImSTgtpzsbIeJNxJpVQ0fdiNF7/ktGHFbQzIFLnNtHh05G0Inij3OWodoaG7st2SdpcU2T92Yp0
ZhP+pHLymt5Lf/inFUt60fnC2XUbQoVboD1THTxGKmjOTV3T7pM58Ig5cgo6EfG0ccbgQ1396+uE
pqJNxZtMD8DcNb23pMycCkDGOlmOmd2dPZjkBtVITNxDKD8dbPkG1vbpntn+M7VljTjKQ+7E3f/H
VXuk2OkYPquhRNwTebvijpfpq/0ga4WTr54LKNxfUsAEz0OEfpza5Nnw0hKi/2/Te0YCeaJXQIVc
SBJhhEGyLScWgvTMVJzG1rDM/RujSIRa3GJ0EPGr0KWBIeYf81YnZM09VGUNo0x6SJ1rPOKOTQx6
GHHmY8Uve/kWLwJyjygjzi6P+mN7Nzns3EuHYpki/eVktXGS3qZlVG0qduAoda7KRD/gFdOMdD9o
kenAb59VxhuxhRCIvH2XrrIYswMFTy6gQoQDtd9MbEeHyFPHAyAs2hMpJwafLwxnc81senU1Ptlt
AWIFRQ0cBzlOq1e38gBq126o6eWWScT6pqfRNE2vEKNvlViP7Rw//xTc7YopuouGnYq3vdpUs0ic
pJvApowZ8+6GrzhFFj5jnImUVy6Oj8Unb4+gazb13AV9aZHh29lgPOnhgKJHa0aoC1r4r1CQKfgi
LQLqQhPDsXTz2fRNtx9R+ML4deYwHQCElIua0/p2PgJnrQSkF5M4HmwdZTdhJci+jEVQ1oeJUkzm
kY1F+cTD1Hq74cLIPw1G39sO5ykHzDalGb0ov1aBIbbkdH7gz1Hpibt+FtLS3FVrEMBSdGLomv3x
YiisXTIG65w1F5b5slWJ/mMffW+QjpBS5qIYHA/WpTLtufqFU6SDykdFlcVZLJdG1udsPQV1RJC2
HbnLXVMSYCAgjEUY/wOruNGhcf030IyMTuhdBoXbQ9Bmp8boiJHdxb2mXTSlCQDkkLlB697zgZzH
s/H0F7M4PcHAgC8D7dsybAmL2bM2ofQUaVxiwLDEJMBjN22Stg34lDQw2dNYAkD+i7M4GCRJSAzw
rlb/sR/kobq9iu23Pk1dz/0QHCy5DbB2HqmLwr/5hHJnhB6TYCO3IWsqldir7e/tAP0sgoTI1xfi
vEmWmXWs+JtHYAZhc3SxMJ74qzwVH1Li6nyS3U1jnP/pTIuv/MQJFdU+t6r0H2Vs4XObemWvMNt8
7OSLTff8Ln/iYbe+QvDxXJtKLyyjR3FPQPd/eLgFEMom+z8gNFIjbo+SIEY9csI84jux/RDyYP1b
8DrmNEpTCtTBkJmKKZRQ5CeMKKop4D5XHg2CXaGaET/ZtO29feOj1hLKRmKVKgD0jQHJnt+0GZA9
f36TROU572X2YaPV891Bacaiuixw4BKGVemLOCtEKPEV3nTUOIqjTEfD+Ui4z0vOKbnGSdxZ6XLm
42zuxQfF75Md9yxuhpSj03Shhp74/QUrVpvTkysPexRBN+wr16rLjk2vP9WlWUxPCc6uPO1HJ2YH
U+Cu0/VxGRldvmYptKQxCs11/RAzA8wCu8NIbqEi5gq92aMjxp31MqYWCvmXzO0GUu10z3KiX4nY
wb876bNOk0qK6AcMDA6kjgRliF+BDPf5AroW/mv2owp50tme3a2w2DSVLLOxwFD2+SU7Q8RwSWyh
PuPSWuxHqFAegtee8/jmpayAW0NWblMqz0wgClxgC/eIYd8PkyQWiUJYSXXQSPE1/P7vaiiYWvzs
5x5ZpZh6sZhhHW4bLQ+eVwqk6zgEpIXQZ3+oxKkURtXFa4HhK+9KPXkGn2XAeSyxrufkIUcq+d5T
Hlj8JAxcahOq5TJ/uLZMY9ejpr7wbtvsAeSpWl/eBVemqycKCjl+GoivEBgCPSxG4KTdDwO0dRBF
EvYoUEbw2Lh6lRDRaAEZ4Km4pedryQ1Haf1V94QYPutnfrfRYOdV5zReVrtLPf/5Yx1sJavmo2Qb
mQLVP6h8hPjdA8Opfaljq5To6gZWHd5jKqQMgkfIC0oCn4bwCmKg9BIZo3mlsl02HxRwEc1qkg6J
VRlnnFGNgRam5QF4BpJ/n5+FGX3O63EgE2irl74Eu/bIByKJKtBPJwNnj3fg5lUJNC0GCmYrW+Yf
R9twAXjOPk0mD/GpEg4yKlxk9uKLyodECLA7gfJ52sJAiY8wqvJYOOg8FH2i6wgzKs7TL9G631az
w8M0EsA4RybIFBVlCesbPjEY4FFYSCC5nhAWZbAvyie/jq/OnbjAwWw4aAok4cHvuomIH0cqpLeF
q9U544bT6mR4XPmjIfOXpRY60lnbjjUN94JWKYNUbgBFkrJYrk4QnycnljK/iusgPqdohgyA9LI4
tdHWMBlR08GdT6RbrNZnk/1aqiwi2QIsza05J2IAMLGdzCbUGsqMMm3YIjvE4FnS91kVwNaMcsKD
AyKYuffaSRJlP07DuP4sgFK02cmeqJSocaM4lLLkwjpijlJs6+5rvtOMEoIUTWWrrNB1/zBBly32
xnbLzr5b8BwabT/pFjYbKymb2CTdC9ldEu/ue0muTMK0yg0GhOaWroOk7KGHvaVgmafCQKCmnfLy
HRqPOS229NYKBuxWWMrmrFUopTTYHv7O+ziYLgYL1TNmqlvsI/DhlwDl9q4Mmtm8dqOmYYdQesXy
LtxhwQU4mj6/+kctazFuksc7GqeMwdlJLl5ptfmZ7JSCo7q2nkxNAh6hkLVtL7cWcUEMQWO3mRDB
MSQLo6FHNEEzWvSIx2+kHgk3a5MaTL1vK68BsQErHN2mXzfpOpYgokloLqMhz5/dB9Qo6eCBhwv5
Nm7/Iz+dNKVBryQqmUEEmQlHsP84OlL/kXtRX4B3xF5D8ShY7etIOukJit8GJtIvTZS0P5JCENge
qw7zxk3bmVAkyqRWITdZbPhukXqaT70Lgkgs5WNx0wt0H8j7AuE6vmHp0xHzuQMjrG8wXPn2YhMs
cNkSHDFwnGEhAYzw4Sk48jFzmb3o5N1ghZPAJzS1grfJh+XvL32rvVf+tWFan4+/agVnM7SNKZDt
tQqV9yvY9jmNN/nabJ5UxKhMDRaUukgm2GgO2LLbz+rc+9jU2ufFthQIXFf1EaeEXb+TW+TiuB9+
x1wHfXTPnnqBH31NdIU4l+H20kiMOUSB10+Uda3u8TZWtTF74whQXdrvjyRT+FWSGW/pDP7WX15s
vki7X4XtUiB9wnruvfNm3HfHwYREOhuF7NPQQIxd9Gxo7nflsdKYo/Gx4y41IR8DcdrrYhukG+R2
7WTCg3UuSz1GJN4+vuoUmokv4MIJAd5e+oa41OnlFUlMe87U+JL6BTzAZVQ2NLaMLGkJhciUgeUK
CooThRp4xl+6sqa7+Us7L3yub/8OWqqun8KymaTuv3yjZVLbtFyZirX2pJZpSzs9bC37GrLrjVnh
hddbNtAc5y7A296+ADk9gm+fIQOSJz2J1hLOBc3TWJSPUOnyglOvq/1dtURTWWX0u1CFhvDG5WPR
TcoxPxe6Hyi/97Yc2Snc37wEfUcPPxZ0Lhu+sMe71O7jZo7hby8gtZF3Qrnh52d8/EkLS3Zr9H9B
AXtMNz6zK8GrB38Ef3eApa6R4fNgIGgOm1hKXya7d19Zn5/0873cZaZk1pCjuJ6tJAPa11UbrGE4
1SsrmfnbHQagEKkM7Yv0VWWGErx/XcHA0To7tvw1QZ993HFRw9N8LibJH7TmuvnbBlqfs+yDYJTG
6AG/DuTrc6yqk2tGWEamNjELMTjpQVuJSy6Kzsbbld6ldnroJNshroDDS7CD7EzLrhKZfP87ALxm
2UI/ycy+PLrFTxzS8wZcaunMiOL7h7fb+uVGnwlp8b547YexPDbisDBBFSwQb12xIZo2vX32Tnsb
QrD/uA4+uvUk+yXW+ReetnhQS4TEB1Ob9sZeMnuSh/YH0LwU/bbjILE4MPMCmWQKHHSNUKFDabCb
+vdgF8dcI91KZePBkzkgqnPtIpY+QaTqL2qqqzVbgy0nLhavhTQYaWg6APH7/isS5EHcqLLnXOXo
sA7UsxVuJiASyuTJ6eYsDvOeJDG7ZymTJIHaRvzHaCsQi9UQ2t0B1hzod40aTmO4Ugg8ZEC25V3z
NxA4xvIQ7uGx3dmudfL77+0yo3NK3stbvD+01nptSYGTWdiVpx1GT4gLe5DyZVq3Yi69b/rPQxQK
WrlUi0SM3EasdMjv9BWekurf2QkeECunb0H9dKhKSwqO4J+vhBMCKuUfQKBnn8meOCpfL2RHwbTj
8bc3yzSh4voVTEvcSSA1BFXUIq3Z5bricOBsaZPkhHw/ZG27OoNK/m4tB646Jux+zVKUfQF77XQ1
2sRGBuIl4jug4T/WiFb1wT/Nzs4XsUpUGJ/XYhgvOUm3gi5mxofIbrBggN4eYB63Jpvd1J1IFQ4h
HiwU9d4DiosaRHpXzqL6neKs7h5U8jBqUBMf39timRccnlG4Fs9JHKEb/NWFZfc90WCYWSpJeVrk
1Kwoe56S7IWuzMzEXW9GaY8fSkhfFRukDmZN/Ym8TBO+jVZdGoE3Kan6K+luqmTC/W8SfpO1AMji
fcl3MVGVy2V9QOlbz873S0q/KZeFAgq5TnSrokL+RbI6iO4iFCeX5fpgSFSbK23DjLNWhysrtW3P
nTYqmJV9+ds4GceTNyVbk14DBkr0X3WSp2RFucSPDpV+npfiupm523Z8HiXef19W6bJuoKTAX5yj
ilV6VBOSAETyA90jCUFkgqOgRqucDJ9j3W9CyrEgoca86orTHuB2FfmdrZJykYIfsHB1A+kVC1vO
EMF0oZgecfwTD/y9Y50iaLqsrunStUR/+nER0mMxaUQMai7lAhD8YkInGZzEZfbX1oMwXVPTXfSH
VfqH10IlSxSfVf2F/km1WbhBPHGuCmqht7Af9WwvBVUL5YgNOo6VE1Hg9N4MBmUg7QUUzt7ADuWb
0rrVov0jR46uZdEL/scnJKabKAi/Cdr+cLbmhAY05jH+LmZtEwdI1eSorMfhBTwNA4LBKn4QYPAK
FZvlNjpRMmr4PA8nOjdztvMtX1vcEDaIf8sJOZcbjR/OmL10izvOZ/43W0o5AarSAWa3UppUi7cH
HGpQtlpL230VB5mgxNYIyBv3Q24tZLqiYJH0OvRPKs4bLQQVanKX9Y9h8xenpQ3d0YRLAn8ylBkP
+19BaEYiWqq8TO4C6BBfjaOJPOdAI93JQaTHznJe6unkyHlVF3BoidtjHdFxmVG//+2i92GZmUrz
+xJI2pKZ8d5IdM+L3w1Y9LBX+yXvRO3R3Kg2hK/dPvXXuCyHcTePLtZpCRtAkWCkkSNfIrovvpe6
Z0Hns7qeMN6+oXQyHOOJYS4rQyFMAZdhO4NjhHWTk7wiofdmYFaAr6SFBpaMBPn21YSsYM0tJT7R
U/Ufpg+0ZHhl6DRHFTFoOezR2m2gQwonHuKjbpJGDLFuzOunSTwXC096/ECcD/zZV4jGc2WByyA0
O1lq5Zy9ApYgUeydjvVDtAu7DB71QxeiEADqHho5hAYTDCGpK83pzSiIBUeQ+bokZflXR3rQ7S3P
ibPDwfYaJGVIRoihiXGlepsoVvytjPXoECWq1G+T6k7bvGZjnhIrVKODlTS53bnynUOIkMZKjiXW
6uWIt/bEaghsYTeAjJTz/LZzh8neaWjzYID377hHKma9/KmfT4qZGTuR5OqVP2SHyg6t6PfLOyfC
wPqf1tUk9N6fnaxakY6iH5O3sxx5MQE93JJ1DWMQE52o5S5qknJI+dYegaeR4ilswG87aR9Hvzan
yn+AsWwt0nA3bpKJrLwcPizeFsfbxx3v0ADLXIYFQdoG15mkXl4Gwr800IBMqownPlYNBYjazdUs
kOPKTRiRTf0B7aPxphcsopcPr3hLaiQHwkKqEEt8Ns3AZrPOg4VgXx4ckPQP7utzDEf3WzWTvjJA
DPB9OU6WFWTQuTVGaFnKkMCszjW3jFeTGikigLk/WZWI53VG5VtdFSi4wNOqJuFmwScxVHJmVXax
7cp195sNjh1ieoNNFefOTuVHbd5YjGhH+n4IOkP2iIxK9svo4KLglVJ9wyeTdlGmHQz80FwN32Cn
/Zo3S3EljUE+mV5nHTcAVQCVDAxcf3sQQN4oHABQgGoi7D9+EM8lf2XPGJzFek5kdRldqPuzxwPz
28RkxbTIBdlMFT3Jxa5iuWe0LV8bIuLF1YAvw8FAf5kL6wyoJ5ISzTXE2IYCQu8tDfyBe30VEZg4
tL8GX/tpqDDl9QboJjqGpGaRINRAGEfLdT4mBofuYLIvUSzdBHNrtpIM/1o9utCzgg1SmchlgQYZ
rIhk+JgAWRfuQDPUyuYV8/1aOzo7MdtuNkJ7YB/Mstcp214UAFC6rpSPdGE2iMi3fMo1AoJV91DM
sfVh4vx5zpmlMfcuGMX6SG6lGK5sTdLfL1PMvtQ4RnZAfjE6feaJfsfZ5KzuBdGqDPpdzHSboXyX
fTFVLsaKxyDRlMcEoMm64mx2mo1I3Xcc09g9M0G3NDqd87aIxOQzRtwmh/3cedjG/241MRgGGgU8
gucsTeZ78z+8u7x4oEDg0U5fVXE0v2nJH5DA3OHhQjdKDS+WOZ4wrI1C7r2IMFEimDXoGFSECdGq
F1EwDnKvH7DiqCHNMs1aUUq+w6Rjz55hFZnDKq1sUtBkd+30ZhW3w6BB+dQmki3yeRP1VF+Lcpcf
BVCf1bOibV3M1fFop9/bn++P8y2mmCz5Te9BpJr+mMW4xjd6oOTVMadOz0JkWS3PhML63WDLQ1QZ
4U+wtBK1p/YQ7f+MsSgLgjoqU6x8Xrou/kczr03t9LzEgbFXF7pw2HF4ZQ99rN1XGmsp97ecAGuq
e2saGsSPOiWB1UPCuzetX0MK61OBpjItJ2N1MdQrvRiR+xBl3TUdVKCi0tB6xPkH9xjZI2uUh9zv
m3UmoB2aseb3vwH+d2bDZNlX2SBxKdzQy2HrWCR630Xne0FZmP5VHg8FGfCzpKbYDdH708FGGVlv
jeAFBpkzdbpoe9uDyOb/6yqnUxaA0KxdyDlds7hsCVGGw+liRvVL/hayvgWxTsFSO8o5QeLe6Wwa
eJUziY6cCJ2X41XvIPeEyN1zPZIW6dJQssk524FhKkE0riuyYV8rg5UEfgKbF+4Juu8gdGwvdMpF
YgrpjgiYUcTIsc9RBgUWLGlFbKRwsZWmGsbfTuaD7GXS2b391Eobe/GbjphXe7EmaSdg1s6Sm89f
YvcOy/FUyYkoXgJzm9iOJdck8055wsZrabVESurWhtiCSz08D3Ou4FxWnvY6ivxwr8YhhNKnMv5E
J3XCJ8jUP7fSK9yra0hWuGTTt4iSeGs9LVqzedTJE7quokOQ9VcvRMdxREU6Uk5t/uBVWv1pDNm/
323cooqN90soW4QesTc5tS8zR7DjPv+M2wgvIQw5QAHRj2PmQYmMQh6GIuHpQDQSp7QpfvtTCeDA
Qd9WYsOrAOm+L6VDdD6yDPgFpaY9b60KocRCsz0HQZDGMLBVZ0nx+VqbLnXLwtkDsBLLyZlb32s3
I93e3yanTK03w3Qidsu81WD218MZ1F3P71VqiNzDVA4U5aDTLOyhr10QY1gtHcXAYTZiPKcZ0Eyu
alVtKCptpZ+PM7hZscZ3YgpIZjflckyH2USuPJM1gMxwpqnnvdScHfaOAKfTgbt3IBLmqUe2eUSb
qXg1v5WB9+joGZgBhHqK5KHpoaCM6iQmRTNlujgsLus3A2SrRJFKQnMUOti9W6YL1tn5abTsBsNq
VJxuFzZDg52N5M0D/xqqkNfn1+8dXo40qaAjweW/NrJQT7mN+4O6IpLlMotHzBIhhZU7uvxUm+8P
b8cd8wq+M7Lk0w6iCI03BkqbXUGFkBuJuVfD/s66NyvtEJ6qH0hY2GTdV5eTHB0QJk++txVKe5/F
rDZI/FZrIv7tQq8qTWkh3PZPKsfVtqsNvoPJlAO1H1QrpuE8rQWTHb+mmmL3jZhOEX1p1vuURxJe
k7RFFao5b5hyuPep9KZK7VfiYmjHrJ84CvOAyWmjCsYYceq6i0k00EovrkQz90yZdcS7KonQmejj
upO5Y4GMzBZnVnlYbm4gf1+a1gRJPojrOCirxm0qlnzPc/osoigTqb7XD/tJnndKZqiMeGklAfhJ
69cAPc6sbS8MnveqVwHlrxJTzv+rHyC5wPsfMozt/k0e4bCYI6ihXXPfwCYPTjTkgH3vy7nRunjT
1PDJ2BFdGVAMyo9SDfs/157KNv+mEICVIGW7IxyH2/O+XTepp2QYevsF6YKULzxWV8t/OIXc1RH7
Kz1ukk0yCdfGXoCEYdWVzik7+yLSZS34WjuHmoakddbBgWcybXSOs7BfQOcPmfIbJMDexb0MDBWF
849DfP3K++vrumckF4uh6TgVUNmqivvx4tfkOtDF3Kn2OZLy+OXqzD46HQYV1Pga+BiltrPF9Mx6
T5EOXGNqthB4mBrwz6WzQKlanKzjEvx2wRmo5wmAKAtU+jdmpRTqKXrxDIaB89peB6LaqK2nFcTz
6dW5IIl4VmPZp3OythMfI/qNYEMt22TmhqdQibMMmJjKpQ8ACPHKPidp0gZgHCeQGnhF6jVzGxj0
WauEbt9mJLt4D+xVi2XHPTdMeQyx7i80qbBB2KPZZAvM4TMqFOUwTPFwe8/fiT9WCWbJN64f1nfJ
oM/k51QarW80AubMgT6iEqcTUi0BaUz20AzoGAmFySdVRtptko5+xKZsQ/P7fYRnWGjKFEiuSNRU
gCknpvJkrgaS631VyjAIyZYFcOxHXpZa+AxkW9w3Iveg5K9KZIIu6K+JqXBf2/8aRO0Tnd2NoxAb
MPiVxPWYzRSNVsLhWej18Aa1eTCNWIFiW3fl91490I+CuCUnLT+Tncf/VJez2+rHnmDvMewIHzFu
LKVA4orBvVK94N0GY/QZtXkvpDz76wzaiJP7OeWEUkadXETS1qvJbI4E055/FfnBkrv3M/t+ZrI1
P66ZpXc7ZkzHu8Oad18L1yXJ52NUamDXITMPpSMhhBrcnFaVF1CELQv0BdKvYS2E03h5zRuI8w6T
l+dsxv4M5362f1oopAGWl2J+SToJTT6qNLasdFyUmbATOAqlI0U6GAPMnArpNmiBSzBqb4z9bEf7
PI7ZwHIbvNg8qlFQNnft1GBVnWAJfYR1x1d5xJvxz7px9GdeBtZtDLDWetmMP21t8LoPFD+c+GJI
eFQiBbJmjbZl57BsPCegx/l9pmU6hyB01YT2rSxjLpzYAKWQfjtSn6Aby3lUhNXqzPqKt7uItbp9
/0K+obSZNRn4XG2jKiOnuotrPe8mQu66T6OOzBMZAV+Nv8xNmpPhEVa4nnyg+Z/YDrLw4F4WGBvO
t4IHh8Vy2pa7Is4zs9DZmjEnWdRM+B8sh+kfZsE7hRZHwFgYUmCCd/Ap0v5k1J1JAXpUsSlVlmQu
tgqabvE7UIRMe+3FmpdlOmHiL0KnslsCTZAa3d1wagnvfDK7v7/6wWXQMlFKG2KaNzL28K1kkto7
a5/mAh86NWO2iAex3D/hrQH/NXzLPkdr8NbeYI2OzRQ9h3xjrnk+ZX1S2ZCfr7lbfvNuoL46pZ9F
pF+sLqhshhYReuPNqdGWhM2BYX0BUu9zXW1tmlX715JaBtKt6NjKxn32yxz0agOWx/w6rPUGrrO7
79DH7TIm2lH3J8eSWoLFWVrbbkLZcXM3J8ajOQJqw0ElRpnl9c7Osr/mg6VRIHfUN3Y+phLaNY0e
tVITEAckLrs33xUIhta8LLoucmaPkmaPx5TF0QrcZtpCSNVVn4XLgGJ233raplLNJRT7ph4JxY8G
h1o3MBjqo5ju+G/9gEdX0+QK15/9LjVkwqAWXQFmqPDIXDkFRatyWfRiMZ5QXaLTyNnxqLb7vWu0
RxNXKY8Pt+HjjLihx/8WPCEkiLK3sCC74sy2YdB9I7mgJ1U6d0j7dNUTgdodoDIBHUqup0XfE9ko
CNLaaLR2In4JIz2o1hwi4xCNw/7WAu7X1Aus0I2xMWTufgs71qsUY3hMYpd+9fjzjgU6bAhQoXaA
gQQm2+fHO1RzM5dEgKUiQUX1aMQ9mUv9ieNA7IbdXV8G6pf5xypfLYkg81tGltdz/osv6B60W++f
0ImImcQORneihwds1tlNuDTSebAZF9GGDne8JriRlF56xsNmiCGuNHjrQF0pOXjG3kohGhW7G8a8
S3m2F5BqNp9mE0EW15bXkWf+Ecrwgc5H65y2tj/rfqPFRvPb0B3ogQOJ0sIBhe40xn6+y4XpvPkZ
12xjP3tU9FrXopX+1nT3zuwEJQGAcBqfj9V7wdxsltBqgwLNlZoU6XNiu4HaHw0pztU9IHz/0WdP
7RFP3WwNNQDBfQf/lvqjf8pidAq48+sS7Zkg3GByLfij5nR+PnVWgXbaaTi3xTBTRkQdzCkEO1ec
m3VuhFRZswXaiCPde3MwPHHimpSMGUJp03a7HHkD+wYpNj0S9GEmMgB0MlBqKANuwQBxvIRHqqp+
O/w/FSTPJVJqNdr3rNNCtrlNh6ufI0NmJN0RKRA/eH0hzNvlbXtYQuL5Crsga1yU2m5Xk2nzEJv+
I4k/DQZzJkZu86rYHxK4T7Oiw/dyfXVP+09/g9vaqGNLFdsKneknLEvAazSmXSJV//ApD4e79olH
+P/i7xlsJcnEp9JJl3qTwi+ZDLcp0o2uc7rFhe/dIXS5NnrnK7vhXQcCNTLYjQ/MQ2yOy3LeKoOU
kvk+Vwhgg5HYgcYT4wYoHcjrvbBcC+qa1LrrurgaiHEUWmIZAps0OAJVMOcdaY1ZNbZjWAsVevZJ
+FQe+k+ZWBpk4pyeF16TNZTQGj4tfjZSkLPP5bHCYJEV6om+aVfTpf4P4xTZd1mKquArgl8n6+Pw
w54yFFKUVTIJjB4QrjFdm6S9XUEcyx6GmzEl5kLu9bL9BRMFXfPnX5I0mogu0TEuRX6plEI5Mq/t
8S4mFKbOn5oEAd+KwV2Tmm8ADsDp8RkOaQEjDCOtlz3n6jdI7K8+A145i9vxRcZ3NkeqTQMMk8RU
kt6RMFG0S2zOj4w1tPouEs9PIJRP0qcorK8FH1gqQ9QrceunXha7jz095Xusualh4mmEb8RXto+1
ntmfgyu3yMAWWGJ9qXS68sqMhtF1yLE6EHnq5KN/PDEMgjIFQEfkm844F6Xno4TBYgkAoUKYvoAe
cV0nEoTCWDjOE2HwRWifICW6m1oZJZREW3dlaW5HXZX2CvJ4CKHxbmJ5yhPoFTj/oyEe5gdd3PYV
zVRLs40fGL6aNJjUKWN1hU5coPJqPwb0+RvkkwMaGAQ2tdM3t2g4eUpUVajKj7mfamNqvi2YUKhU
GOj1kUsPf8QMW5h4VODURJBYFaTuwRlprwFuUszlen0FaUgwqe66FTW9SsIZS3sbvZA39GskdWnK
RXg7/TusbusPCh/0Adn74RhUYqtzEHxGGwEjX7ISBk3ueuCOd0RNCIL8b3MSUOv7epMuOM59zQ1d
FxF6zw+leFId8mndD+nWC0hXnt4SI3mLU0+0qtU826NXbQ87FU4GN0vmkqHgrYEuyZf0vyyVYVJN
JBVtKDXkUjA3uznvogCK31kVqwPsa2TdFdgRgYQZBMMa4Iz/lVgc7wRPLAFN7+oTox3RVMd7Yd79
dScm0XSVGALWin1QOS8gEv5nOLzDzaEHJQLCOowADJe249s4KnAmLCSMCQh65muPudjN1hFcNAKK
kuslZ/VYCH7UONWQ11TmboRrsm0wnayIluxxNPbILHk4kuuhYX8UhdEIwFd22BpGtv6fUZnLSLUg
//zlWvUXoVnMkQv5QJLCjQ+dSUmQFVCvm21hc6j4hDXdI9wNhQ8YGO7H/HfqOX9bx2Zb6iX6keIF
WO8/G7t34hU9bgUMoRkWBywYlWaZTWGmjRvdjpRuKpp+7iNpzhHbYnzsWm0sNkqvX6JAQhTsFHgv
azsQps8tU+zK8Juck/whKewDXpUIy7qM9aSbDxu/cnJtWIxFbLshEv4DJD8QgZ3t6/AdMZJP2Qa5
gDPbS7KxauUpa9G4C+LmiQ9Nq269SZVvNxQjXfFkfhfsnvwRJXw6cSoPma/q7GAQXmMi0OXpQlbD
+CKbSbQvWBPnSHNPeeQ0oVlSrZ9oty3vwuIfTG5w/hv5TibRZE0NNB8BjF4+ut5z1fs4iknwfFCu
Y8MQWLrxAuHXA1na72lH+tJRyytX3aTLCQE/c4hXryQqgw1mhgNIyjgeW8F4WEyXAYoEGyTjnfHR
QWRMTxl1rRxbGcGLn2t50aKorecLY9nzolXpB6CU8UE/Hlp9DU8pVAuNyGb/0t9tdDcqT5ZMvUXy
2t1GzUd/yw21VdzTvgnnuyiK6qmT1eoEkh82jacNcxhwkwifUsMvMq3CsSdNUHdfNpXC9K4QF7Hz
B+1UWMgJsi6+6mhFAAmFDMnBCbZKVCh4tRVYlUz5cQ2IFkavZPFzh8R+M0d5iAvxgon51SvxAlJI
ZaD0ZC5lOEGim2xbwzkdEGumaAsLziI4p6rcNsfvuHa++AkwOV4xfeeqYaJHeB2zYCSVfENqEOJE
KSQVUhBJUsq9CuFCHQiiz5fNBb8YFBiHnzJdYl0vdLBpcxEGInh1a9aF8UpJbYH6FSCK30M+QDjC
UIKcUFZ4agf5erS7HnlHPr0AHS4V4r4UNpFsgg9/MrMsEVQzY4cApuGE8TN0h5sgPwVpBrmpSvjk
u4gMMWuBDLndKif6D4/60zmwErJ2dhqEx1urCa51h3t7xFGCGOJMZhQgf9JIc15WoFXf/1xZUvBl
5PD9iVHxSxIFceJWCMwYMmULazTtFNjO+5I+Km1QfARYIquhrDhJ3CeW0Yio6dgVRq04j8WCA8LD
8eG4EhhhWg6L0ucdCN814cURTxZkK/K49yhNAwHTTJWplsezuiEjrHlKB76Mgk9xIVq8UTyZxTRD
4YNNhPaGWlQkdGTPhaGY2Jeh5qVMza7uCsXMZ2IDc+tXZm4YWlq9P8jgOLmQ0BK1qeFrhDyRzoE8
yEQ8bOwHf1iRqd1mtUicD5b8P2gtr1yOnt5Mf3P8IkfFtvx/aBRmTMbIDUUmMtZ/CedRl/EipzUY
FwOu+zD5b1xaf2vjb53UqltshNs7ygtQ7Wng/ZwmtAXDhzhfvhSBFiVPY6fMtQ6MvbHbGgzL8MTW
M7WOEoMSowXxnQLBBHvsGB3n3sE7pxU3TQE36TaRPNVwnNLdPyKvBtDh4ubp6mOl4AwBZ5zOIlx5
sepR5pX07Bke7HngO+nxzveI4iVplZEKU6dmFbwUyw4DZxAJyU/dglxo2nVfLyE1pH2GzMomOlCS
czJju9zH4Krgs8CnrRJvcBRib8hvwPqAFNj1vNbMWFRmAtgHOaD1X/hWlVV93ur/JzBbfOoFHWE8
iU+uvaiXwggoWHTHTyVrEyvJktzYRqkkkGYRb4W3c2SDdLA5EcJRYx5nP7dcTB64BZm2Gy+G4QGo
TtNvN6nETD4cNOOLu8vJGH1WNjX7MUACbC9pcYTOmmiP0f94D4G7xSixBDU/I0h3Vf6lrfDuJsnc
I1BjLZ5Yh1t0yZRL9Qwz1d2phqKLWK9WqsyGk+7RZFF/Cz8YhFEYhMTrwI1Ouaofzm/9TczoKCDL
m1A8+VtWtXyIZebeHqy46ukqlaB0qoPhJSsuyD8fmTN35DNtte0A8uhrWxzjESPEnmS7/P5w/cWI
6SLzfGlMvmo9M8CxRPQcCzGRCojpusQDoxFg36PyIHs1JR62bIBAuakuce1k4481aiVnMjRuKlRU
iik1R06dHpzT12da3Rn//mxJ4Zbof9rUHIKg5S5alhzPTJO5LHNKee++jX81QnV3aXz2tFeAlQax
wq+he4Sm1Gs6KGnhR0UPybeUJyCjfZNlwh8zQOvshlxhdvoRMFH8ue3xZodC+2MfmHOJaVYik8X7
ELtVL/JfFYze/9q28JYO9ZOIYpPVrLChbRqN6hP0qWWPGjCaLOjsFLVL/guELiQb0oqbdagUG1Wu
uxWMKnACcIsByQvv8U5prYYQRW+nIb/AkgFovCU6ucuT/aPJkKZEuAOK/gq824hPtS/gu0z5Z1Ix
S+mrkOloXpu6162rfRODKt4M3xXC1d7JutlzHbWhr/MIQcxB50q5Moc5reovjKSFfvUeHovEak/9
jnXfeChoec/UxXQ7QDgNLjltRzL4VorN/kl5qcGb6+NaPgOOS43htk3SGJ93a3qQZlrlzhw7QLtx
KjmMZquPOjiZBbvUq6HVALCaiE2eTJ7zGLzOBlPXvUjaxSVJwkw8swWRiFuB2LaDm/rQxyRDzNWT
UPxePgKZBh1BRytxZw1EwqDtfuWOPXkpBopZtVXmYr0v/a98g5TbPACD1gRT8gBqcZZaGyFlDw3n
9IxpgW3A+7UedoAX8bO3xGEauoz4vwJxeUn8aBvSgmrqGhC1zCAZTmNB1jMyLYGOmCpBTIgGanvO
ehNJ57EXpFBeokAWH7RQPuc51quzp9oMAq1j7x0ohx302xSqYsKfJAxaU8eRFOQBjQJ3y6vH588m
6UI3IVPEAa54R2ojA2mKp7QLuCACVtw/hoS6cewyfwevdjaxT837huTFucF3w4dGMbFHjMgBLQRd
Jg4pnGZ6wrjP9FQlaeh+W29mSGgd2C/hDop3HBC8fihgMx4IHeUNfv3OGY8NVnsv8n6BxeqVjOtx
7kZGrP6NfNgaQ44YoThJnKZGRRYahaVXTM64+29tgfod+ZljINqC1peWZIpl68Ze/2vh7JOIFTSj
MVmM/dBBZFRlFFkHMUzZ7HhhiqV7jDG3nrJW3E1gQD/8u91AlBN/GO6yd6KtG8d/GsoGlSWCB1Iw
nk6fKN4FI0GHeSgz1IO2sNSKCnCRydoeM2ojVdDBslacBpvhlsR3WEqX1kjMx0gC0ZUrNnTg4Ybu
kJmXbIV7HTCNX6fXXKv3yUXmomX2KzcQXSRu3hILXTmTD4+st5ZshYUniH63HMJ/dfrHOjT4Bfjo
M1c1NFrpp9quyTgA0G2OgtXQKX78NbuyslF60Wz0her267OuDSGTXfPThy+kK/DvCdRyfIEZyw2b
tucUwlMwYFbVz7htUJUsQz207TPQmZcBlhDCjDoUcHM3/nuRIrra2IVzDWAaL9B2Li7/zlPeOocy
dIeLuGp7PtDLhfQbKYRhND0UefCgsul8og+AxysS+wKW9j7G04KAPwDmfYQ/O+TxbGcdL9O+myvd
qXW2u8nmve04fNqA6ejoniVzBBNAlik8msmujNa21cfmyZQ6Nds/VjAALKpThAlUdBiDM6F1zuIA
C9E35JMGODQh8tj/Cv4HAopPE0EntFwZPkZoAn+sBz2gBHIRn1BVhL8MbuzUW2kD4qvM+tYnbp83
TAyFEUdQxnwWGoSioJ9Et562odKW3iIKwAwZKHNX7cAIHB4/AX+u5raYD/PjaQ7viVR0Fv7Jughy
eZejxLzRjwvcvkS73pYwkmZWB5kn66ZQ8NTeGSqrXlvd+uSLHPbc+af9zwVrSR66GI/ZiqhrLEA7
vUnesiwRkDY5kOKVvQ1WimzgV3UUDMIXUbdGNXSAMrecf8EG97eR+xG24d0GtTu6oHiLyV0/rmgn
exypGoluQWaa6obP0C4SUvSb3f/VMPKYpihx0dZzpXBHYgWCnOJf3J4is9ONdfmputmlv2/yZx/s
ZFDHKVcVAkJv4RRqczYrUGsVpUJShRiV/QJ9j18qB3qdc5gbJywaWjMgLMcgFVHfxSf3xbqJQAIA
cgn+v/0tIzT5dT7OIM7586WD8QH2rfsfdPOjnfjkGUE8mydfFDTvlTf783dke4Gq3SNc1XX+z38a
he4D+5WVenck4qXkklfcAsnTIlOZuIUJ6E+ulrpZGSEt+XsXtuv5didkimm9qrTycvWCqqSQnSF7
aRG4QtM9vGT9N/TtzBscT94giQ2UDh7Dt0mF3vBjuX/dwmTvl47JSz+Q7P8I3HY0Bwn82Pwg5hF4
SccO8GGiDbfTLM6/HXXb+BhYuJPQMrWA78LIcG9io92gdStfJRikUNAbIcmlyL6y3Gr+PHZdyFGf
CXiBmF9Bvss3MOMMGlewpO++43pyZixA8cS+rlkO89sKAOAcaCkho7DDmdcfT5+OnXSXohwHwh8w
5zGYHdtiDn9o5znPtx4XbHcQKuoFOw82+2W5Nq1RrqHuC2+baguynYhODclSvhzPMLR9XOYrBS0Y
ZWb0aTE5W4Q1DnC/fBhdWzRTVeqc0WiINbiYOYoLjqxUQ2ZZ9DP/u+WIcV5sQlachMaXeO0egg/F
LCj1qhsb3QqkVVpNu+oonXo4fhMkCBFU2SYF2IgupyNYIIfW3Q84TMYwpnpi/ERNVuN9//vX74tf
w7uyy2zHSzEOBWeXCe7Idji77ZzjxsQOpV7GvoYeMLyXNza2hoelx5SYkxOdZybwaDGoSin/V6sr
wR5FZVQNnhJG9YNB2xCvF90tujYL8wWkOeRD94FGq6R9iOBSSOMK/Sdwf5a/3gJNA0D2vYhFQkFb
CEVnQuLv+tnOVzraF+lZHZVc778+8aPbSIsOEYKNzdZXrd8HqwrUbi3sej5Ma7HFzvAJKFcimm2f
Ueb5azOi2amYvBKv+2uWgb02ju0KxXH5qJY1e6Yl/QytAW4jUwPt2DqbjkJQTelQAd/pqDhGNRPe
8AkfCsDXamcViw/c4yw4D/RpaX3iWspbsHcGAyllYrqglsIN2NhOXUwq2BVckXVwrg7fm7lqUIDo
051fX6iBtWos4h5EjyvtSz3fdyoskSwgP5LMoLh8eHSfQ10QtwFezKo+pel7Y191C7oiaCz768bb
ytPMte9jP0NY/k/Iu9r0ag4YZXWTh17JohRdqt4R4FUcbYJyuhQUyXfRP2MwdU6BRAd6KTAHRENP
BvhgS02KrlyIUrmitvY5e9Y6wCNZBoYAx7emhqHIOeFM1VQAVn1IWo5nCYdkELy88ARAUZV7fmz3
30cYpPSaQl0sljZbnuVC94sCb9vyUwJDIHJTQ7w8hW7VIYuNPzsWp5bdoSMMlxnKw9Mtro7GsBGn
rHyKvpu2TM3abvMimmtSQ6KHcPzPXtNrnJ9Oe8kBo7EI21ApegfUdWQ3MAXzqechlK+HlunYORKI
agUyiX2vMNXevH2aFWkFXJK2uadsqOeet1RvgXElIZMskKR+uRlCihM4fIaiU/FpekgxCxlWxXDF
tuMY+8FJlzUOyqa//KXE7dMI2RCpNY4yIvkDFqBQTLYqKXjsT+qCkyoeagLtVRSd/9D5ysWVP+WM
dETpMRUeEo2C3Ra3NEyblG8YarCXIC0NnVj0CPo+UtrA0eHL2rNQ8BOIsEWpN0oQ+hDcVEZl33BY
mz3paagra+xlMuejTVSC0ob1xhwLSTAON/htXutYxAlSPY9VmmDFdvEhlI575UI3IUrW/Tj+gK7T
/rmmUnBAZ7p8XGgHcYmmL7+2ix+0MQpmXvY+FTzxvad9qZFgWoRXvt9N6fNWLJq0ZR1lBN/vmHvr
t5dlwpqlTW8U73rcXWkm9QF14vyCipXVEEUYgP56W4oQs7fcXs4hMPGKYPatYOAIda5xJ3VX1CNG
y8zKPx+2b4MDiYo5nM5hVpRoGl0Gi+LBWoM7FoYpmEJhy4ihpDbFvb5YXO3qMomvqT6hSLhcSIti
Vq+LGLzfK/UKi1jcL06zxVTkMw8otieHpOHk/kyFoS7UyOX3QoUiypMSFhVLWXvpmjb0axwUj8vO
CxvO912oE0PhLZaAReieQPc+uNamu5jk8FHIeenFMImplMwl+QUKw9P+sRiiuwCd7UwqHuJsF4CV
Y6SwPfzY7dyNNy+HUywp+dMw08+1vcMMfQD2NG1hQDsLEEHSiQrMuViKQgZZWw1EPxQX2OzJX/Gn
OA4KpUxk9j30pbTqXkWcglRvSy0q3wCu9Kvhcd4fsUKMehzLQBo7/SnVFhL38ewtQLTG+C6hX7Qw
WEJ+NSeC5cZjsnvkmqRWwJPO+3sKZbZmcxxkepBrxfNt3VXk7obGVKK04P3hwzenrqIwrD1hu5h3
ZWyraYi9vrh+wEySp6vS5Yh4gPWc5A+v8rUdzifYX1XqNbn6sjA/8NonvsNef2qyCQpmxGKQzisQ
HrhQa0AW0C+FFRUi+t2uRhDVYBJ3XYYLTuH2dvOmyGTo3SDfUUTR7r3jpJuY2PboOcV/2GPKfS3E
9iIIEM3mVeeeAOIWQxPcWQzGFxsEf1ijdwnQ15YPfts+/p4sH5JM6KqAuAn5L2+EuZE6koJg4YB2
h5E7EVZDHa+HiPmKrXqOzYcCTUuXmKLmO8gYIYisr4PTY0cY3PN8qSHUjlvBPWhbxfXGh26ZPFp5
FOpC1AmLH6NUvrMmKlkoYZRqBpwbf49vvelxQJjMlJv6kkvkl0iYVczpZg+tEN1/COGerhTG0EHg
oi9Yxhr0cSLiySPQffihx8WftBZeJ2MOJ765AIHNVE3ABYweXLUaw9rEgdxg2Mn30BelfbmIVfFD
Tddg3yXUqYBgQp/1tM0xXbl/tfcFgcVxpY2qrf3zWYmvTk5ZsxLfp+gmqTPni3UQSeoG5cisMauG
70SFZry7+NRddHHpX5H33jAWa1lsz45gVJLciQrjSH0ohU4yy42OJZ9dNrCRCqTTO3mgtJ5xMAmw
nYP9quCwV23ZlNFMUDYQCIXhADkzg3AQbuyFus9kkKlq5um8ir1npzqPfobKrQKao7OlfLEopbmZ
rukk5+FbdQ1n2jkPgmt0b0W06ncGIz+SHnumD/g2gZLH+38vjmkewtxOWySYvjFa5Uv2vsuxPFu1
mdJCPmL8gTuTmuEr9FHxdFmeKqW3r1TctwmzWkYVjsJHDlXRZW6XjdJ1Axy5x52kuJJ9UlkxDaus
3I5gwbvnWpHxJOW+f0bUIZJIWbwC78XNWGAiDimVVVMdNfe003yDVHQREZmizgSjDf27p0LakCLt
O/qUWNgbggOPwDgREc1cCR4OUgDZPzbCOMBZfXJlaJF9+ZICtlKK0ECsjf9E1Zwmgj9tOyTQ1wsB
aJpZEsrqb5VEnrv5h/dKKAU8GWnky+1s68oX+5Q4l81Li5/fdxQnUOi8C7A7UilBjmhibHqIMg5F
dOT0HYzVs1x39pgoV34aUI1XvyssGGhLVjTSQyE4TQe/Y7wjjv5pPvWoq9pWCn6q0rRyvD7mKWVn
jVMCBaYbUy77UD5WcHpQIRZerE5Clr05zoxXc4aFtnVM/1F4SgB+ZAqEcdPdr3y0uN4EEEM3H1HR
Tp12rjsdKb0tslxJvTSK0/gMVi1yiB5FxKxWMHer2pvjE37pK07LXjLpECAvoyiHatPgdGrnb99q
ReE0PtPTOeHLWuvCbGHH4FGo+jhoIDKgWSYyzU2WWqxz8yaLNq0oJwn/flMhs/28wkIAgIoHoIAc
gdBmg8WcfV5zkHW8uCqep4gXEfj1KXn726OZg6nta+yGAvd2knqed4JZf8bmgzTfBW4+69mTW3D9
LnB5gnSzr/MvJPqd54iG61ffLX3tXfQcyxu9TMU3MIidqf+eB6G3UomffhPFv8ZWXvo8EBWQ2L1p
uLKpQM/Y1TfAqnWHw3o7cUY2p7rUYIs3ls5uD+Ceu4EfWpOqGX2tyU8CnRhF2+gfiC3dcDDqLpgI
pQ6UWeL8R+qB/UioRqk+rW2bDq54yc/uLpG4jmAWbqOQDEEh7dx/Q1UYE/lsvGrLP9/UWsYDhKMl
NFwDbfY9kEnsi/c63m4Hqv8A8Sm0tXkEoSCwkhyKRC+LH3TykPF/bmALA0HArXDz7ohi+PB95k+G
JfXi9sF6bMgw9Z83fuspdyahO/vxO2Lta9W38nNjLxFYXm+oR3kUX3A4D+7tguAxxd4uayZljyxZ
gSqilEw5CTwJn1uTCYMooPJmMRBFP/dGh4kzWdzXiC4RGwIkF1aeTWnfHTCzgmH5FUidcm9yN4s+
NGpOq/VNd4oFg2QIldxDcXl7qzrucg6GYrZ+RbQOHY/BjgnCSL+244RWfKY+uC4PkwMAuQDFJwUJ
EqxOJ8tlmWF7UETjQ/ZJgiAiPKk9toMqc7tBaJI1W/oNfbHgzAANdjNR3eJ7kOxxg1wxL0EwidgL
r4LoMfcDfNE+Mqsz4ayhuyNodLxA00D9RlsGwijiFHqz3thgIl5vqSllR9rJBwvxknxsTsl1ZY46
VLlJyNMW/wRG4soUsoxm8Me0PAvYTNOFrNJKT5FAxYH6VuIUw0E7tNCmwJfBeS2SBjwrCaUmCob6
eGbKK6lxJGnjx1yEWxgxvpFNhI65oO6OIM55R5UiN3EKzkJ3xJQiRkvAWO/8i+1v6jewnIPaNyaz
cROdymlvL9dP04hxOcHVZQ2fPos/B9KTqU1nReDzOSQ4Wku+9izIQ5D0rX1i36CrIFek0OWpVfV8
bSV1WnwmW3KAMCT9yco/FjTaeJMLWCS9+4yocT5m8G8JlKKGYDfagdW2FOmYV+SD82WdpwiVSntl
aI2GU0MfptI55JykY2OIUo/3bJbLQZLLOSylJ1nubXy7tWoJBNg6iNcd6E4jUhZbCwAHt1N1iZnQ
SmSA6OaH+uDj4jPaVrPvcdnart94aFBkXmyYMNodZFv7uryhih0Wz0/Y5n1jggdjxZD98WaqFaz/
hVZdVy2irvQXEuUXNtJ3l3z7x8zusBjX7ZUQ2D0xURvU/kw7vlGPJujDdrfYCjaPycyY7GquW3BR
3cJ8qEJpN9TGIknfgrfjCX5BSQftkTAuDx7yMxBaUrJJBIyECrwuF2zaOsYWE7cVs6/4iuW6fhjW
2uGk3OBdjFQVccwXmuuRXqLSwBywS9jr6vJEBnKUgLQ1Bk+e5tru4JkF2Nqvc/T0tKGiiLkDopK5
kYT2fE64bEoruBXyz5gyUBcsBr166DYmSdN9WEACQa69s8NJcNzKFkARwz2XaftnaHCZl2d16pua
8is3xFDeveNtq5rKMvTmr4ZRV5WIy2E0QbOQFezpXjAw+R+PaK0tU8FpqqSfwd9F7ho/zuabT4Qd
2KKCOdpCzMjYJYS1Q5SdkDoSWmBrTDomJ3R4mnAP6Phz3Ra2uIvjtEV62/ivJtwKdO6KSXgBdjbE
A+ajuZXqhrwbyrtP1/rSOBRWQ7O0VRkQ1L+4N58gyBKEhw0ogpmYQ+RNS3ixHEVIZqlGF3E1Ec8+
Ngndgls39TEKzbEdVnxZRFJTibJCICD0pXriuUv7zesbyYjerzwntCZWQcc5AndiqR6iKNZzozcE
8JgMui7XDmlY2fLOarnTFpk15ShnQ5qOj9lM8QGxw3NxGQPzePPGyRDNNfefEHrOFuJynymvoKmt
9OuQdxDUNeXcnIX3QBgaL79Opgysp91rYsax4x2UoQFN9OwCMhg2mHf/XzDt0BdWUyQKEENVdGSL
dRw98Ss8qJ0+u0PZG/jEWGnPNJeQwO8L3uGLbAHFJUS2koid7ZfFdu67Kllr2DcrROlhqw/iGE0D
/YUCl/8OB7aXQALmpUoupDERXOddndjjSeBGUEjd+v1sMWQPIEpugOwTc4DBvK18MTTUkLI/B07i
J7C5BLC5LomRm0wODPgMAypVrpwKq28nTRoE8CEtPFBWNw5CyDEAFKqiuRJwKf23uswLecczos7y
nWpZEFjUUJfXr1/zYgHZq0CIc+hwVcY35DHCV1TC1pB5RMHZrb5Z5g/yk+RcyMIphMBsxDDIXWRz
2gKA9ZbtbX4MShuCLJ7z05QdV5SwBNCu9KqH5jTfYCrOlI8+ifxuQmWJHMRbVjIMOg7kGE801WEd
LRdFHIikHQZ5ChEkTi/fn99Ho4BbhKsiRTxIJ8zqDbUtHWeJcMAanvmcun2pH6y6J+NNqqSxyOlT
l/kO0RVyajECSMjL5B+xnsi91kpkWn+FaMSJNxYYY2MyM7ry5q4o7GI3beS7andoAkG4fMjY/bBJ
wRU8RJAlrJVVxRGh/rQDLoqOqFDs99qXqpKWWcshBktIt4sNa/PpfJVnfCa0LK8Id/WUHfc7dcBu
J96IXQdiC69LIsdHkBlKQh9KW48trf4HuzD7Z2n+zxN0C8R/C7KVznPZ9bBRPaNwBsv0OJdZApIh
kgLbZ3zakLjXymBxutJCepEXrhSrbLj0nYxFMhhXSjPg2Rk856+iPy3MuBpcjS8cR5lT007sa99a
rUWDAuAkHzDKF1I7lUNwASZFNbaXlUh2cPJKRg8SHdGlFFjRKxU5dNxeE7ZoN6fqaZJ8IL85A+Ad
qoDINS7GlKz/TqF9mi1m1mCGImeJ0ogqwaxLXkqXC325QV4OARLsZ6ALZPEsIYQw3/s8zEbCHkOh
om0E4hoT5e8iHrnv4Exu2/ovTDLybttM0vE//MJ90j4Uie3K5OMxXu0FkFRHNb9bFMrK2HNKkYnp
8/iYecGmeSk0mCMTO/tnYWWLRVle8uT7psYghOTWg8EDmKEg46PFKUmGK0j9SY6BYbrX5X3oi8hZ
9XFPwwVl10PedcbIzfwtAt5UsFHqx5GnyNZe6NBz3SW7mFIIkXri2WZkDZTLsFXUHQkk2YQAW8/y
gbqS7Cs4TyrDBIKaJa8/OHxsx6ACIU7E3y4PSI0rIxWc5RiBNLyB9EQRatILeBGjqIzBqEhWOFRI
f3CYYPNdKY8vClKuQrNQOFVZ354iRANZpNRZ8sEIfmMrpyfCO4aHz6GtvgG8zpzJpYA36+LQvop9
Dh5ZqMTnDScy8WdgDlV0DQLYArrNKkFZhq0KB1+3r5638hA+pJv4DTL+1L5zNXTJRwnvw02Iqs6n
k0rhaPu8S/62kTRn1SuBB3KmT26ASven3751LyGNFOREfm/0rD+uguQONcWwKnujxCUA5fpXagAM
YluMxXTuOq5Yt13Uk2Iu2hfY5LS6dPrIsZTtB9sLIPdVgPzA8DjP5MbCHQEuoszQp+cBFOv4lpyG
iW3/NSaXEHYpUGfiAub8RRLab6w8OMFPCZjK8Gf9rDvaDoBjAiWdtlyAOb5q4hHTr9gCjAsXt7OJ
4/ttUk5H02OhRc7mkEpwWKj/WOS6zOXb4//Ec9ll284kYZzOzuVDzZ5yhlXZp6V0SaykA6WjgxLQ
2WAWApR3mNLlrlZxQ9YqOBHg6yTh0lcXIMJ65p/DyA4Ph3MZsW6/YTsTuJPn6bfWJ3bvApRpIEBz
cDv/i/803kB9MzNHDfHwOZdCm9aHNqsBEcLFw9lUyoXCyIrAJwiy2rhnankOfYhaoH8BTVRlx1Xj
PklDYb1vszhuDZW4A10Fb6C9b1jO2Vlu1uFS9qtx1j+EuSLa/o58daJ2IYlcfiBKCWxQBGN9wRTR
r4kjqNjq+siUeDwpjpXLIdRKXnAiXXgVyV5IBEE1EAGIVHNdUQBs+vFVZtEPpMqpi9u2Ywgwe37P
LG/NNsyzUhhB1x3jRjCGy8VUZ/XcHLGx6aIUtY/gks2epvu4eKPW0BKc5aF4hXq6LAe+kaFaYnLY
tnrALH77Jw7ppC3aUtKGD02A3AO0slsu0R5nplT99ehshrTsguC3DaTkRRSVfFi50jxkDpy2mHd9
M9ALT1bz9G5L3k65XceiZw6vt4RhThBgqiIJRl9zAycu2+qcwVDNKjY7M9/jQeB6GTv/WsBUZd2j
sX/4GSaUR884S3IgtZfnnRtNfRx7UkqVglhpDQWgBgPmq0CmEH4W8uHDkG9L+Qt3n2Bgb2QUV+8h
j29+I+uMKZzPv/ndZneu63G9pxcBSdXBK9++xdXfXK8tT1KJgYmWW3kqm6vRtNTFAqcp2+pr7Iro
lqZj6v/zuBoKIA+Jz/8hQF6LyHdcUIshN+rdCP1JKG1lgYCmfwd5jki8FQjuut6YFo8xzmNwQ7j9
DICoKFFGcW/cEz3caz/zc6m9Mlfx3lHLR9Q1Fp7zGFiKwKDrBh1rEJDvbIWHZJzLb7A+X4TkzQpW
2QMPUCjibx+vcIfUcjcXwWuGNqZ56T+cndFvg5IFBaHrP1TSoMoiP9xKJhxWARyqiTZsTAY/o25K
wpcZAuCvmwI+os9rlir4lLpKDEda8v3LvhzS0dafgUWGtqU0BgvPgjubZ7MBZ+nNfWQinTl95yUO
peBVRmzmWtBKzZHYf3T2CnV9hCUpE7X2PHoH2seskgqpsChgA8RiFfc8MPgQsL1Idl/TnRfFJXBq
Ej/TI86vy8ZhqdxPDF8BkzsxmqVkUM4hlX27DN70PbemUjtW10zlawoRpGecSAJGTE6xHhALSHp5
UnMqcrGNQJMA5eKvDULkvlJd7H2jQSieHnnCRbEa/GiaMCsmIduofeweqJihmOtGGFDqi0PvOcHs
9RxgMkqPa3TEQmf6VvFk8ENhQVucVgtOXOUYpO3T18YPGDAz50SyWHMm0EuJeVCh401rC8h3OGre
+eOQUeE9PtqmQmJchSRV1/O/S/Bsa/Vy2QKcTbe6Sqtd8QSskIlW0hJoGN99bWDDh3XuOVojwobJ
5ptN66KDCgSGZxSvBoYjj3u8QjavigZ9z6dIzZA2OkQZ3RESBvFZ1lX4Ef95xygcVrDR0CPReIXG
pGrqdl9PDIDO7KVjX08OuclGkwEKgTLfuMeknrK8afkUGP9/w9K+2gU3Ccc+Xb4a8V+Itv9Ayl2i
cywMHe/MVZNzwtFowrgO7wKUjXkjSlbG3/j+UKn2xP5DgE+MostL/Z26WRSA9OfJOXLt2Ecn3vBp
xWdcf0eV7+diifovjgLmwZJ4xBtjSb5i1wxx24koJPBPbWkwlqO45HYkuwU2FYKdxMrSkWEfqG6l
S0Ey1DOujRjG4fECllYMy+vKykm51iUfqiLYb9/prG/cYw7jl/gDavs7gl71qt5hhTQV23twuRso
zs54pEbb1uY0dq0jX5FceU78DS4GZGSKHLUYOW5qvy4lkOz4YTlFZX0bHzg/VQvpUUWZKQn1yYfI
b1rx7LKZHalyvBL948SnRZZJwdjyudtHXZNYZTgrQ9ys5LHacajDi4cPDJKu4q+2QMWzuNIqaXzc
s3JGoyz2RsDbUa+tfC4cbkaPNhfZcIXjyy8l0b+NTKZUvAA3WfGbROKx2oLDMfiQhSUpemsQwNhw
5WSpRT6sjnc4uRRamzTptzCJ5Hh26TqM0W0DBps6XiTLL53RFNTJVh362Z9ZkadXlzqw2meEUASg
mXWwLcQJems5sOSpj8ejwITUjbpCPI0Mnyiy4lPo3mmqej3dwtiI1hStHVMcGNg4d/CNsfT9ftMo
C+BiLevC0wRawEF9OWcxoOvlzscuJcwesYxR6VLSar56kNdD/9ZWGojL2QDYUX9BT/PhiS4/wTEn
TbLWlc5bFai9mZT6w0Jk/+7C8aLl4eectT1kY3PUqdrkTIUe7lOt4qt6cZ2T4I3GdjqqSLBqrG2L
R0DseJx+grTWop69y8wTcXFY+/glxL+F32d8HyHie/cB4K9M+dVKlZ9OA/Cb9WLwpMc6sC/997DN
Z0XuRJJ5PEbvcJx5h5zZebtEoXjN2bRS2EzSVEAJohdwPX6ulGkBkSSNCb367+CeS4Ksy4FnYgeT
CrPWyeLR9cG8aDdC1/Av+P6pPV0sciafoWwg668wdUMEFIL2N7Q2fvzfRQ8g+ANtXRtva1Nd8SA4
o+vv7tOVcDIGDaTYuUFsDM7deol+fVzVeMywTzs92KzXHnS4yA7nuc5CFfrmVJT+E1vPJMyFbnwJ
Pk47rE7iEW8VGHwCf+Hy99JdtXNFkXfWgi/jNz7Ia1rPUm3zO+FGIv0tlUqBFXvDHxuMrCVWHo2K
GTWbmbp/QMX0Vmc4m5mCRE4lKBMRFJoIC5jvfbKclC9vUWoAJIEtp1Hf6pIiINjqERcPDFjDdS6q
aXokiajMjKkEjD5JAJsOzsrCUHhRlzP9uz5eXpYXtn3PpcMDqkzx9abu137DNZ/IIt/OEYOQvW46
0jofsZWhRdrhPQOZ+YFQITSYu35HGLDXL+tEO6ZT8sLP9ZlO+tLHYZVRJVIJbLORi3E1celFTl1O
f9a9t3Psu/Mjbdh19TKIFVFYKtl11hZrpcBjEy30n2cXWLcnC9yHVcUoB5/PCXnVcxlqcRUaCl/M
iJFqBsm8EEJUJRdQUAJsA4GudLYI9f7RfDxbwNMRrxOs2p2b20mPKuio3r7uIaJu2RrRMNyZaju9
KpXzFq3HPP2HJ46Oock+6zW8Iyo1rhvHpYxOAw30BNk5nKDXQPZVmxf4l2SP3/k+LHDEk9w2F5Yb
+keZNyEJiUoHL32NZ3PqvHEMq7yGTTxo4w8onUTI2lGCWFtISOuOseCtMdhLFMImKQi3RY09CQct
I/uj9n9dw2mzfASzUxal42fDfc1XaYiN8fuQmIGIGRrOVVQXMH3B4DSu/5h/UPWMwTlJgTAmm0rM
KX2Lcdg6r10qbNZDlPCPWANkTeZuaKGxHXxwP5LW1EUKKlW1IsVbj/DJxN7PgTseDYIm/nnFXD25
5LWkUOJUMg2GIii43M2QhYKFWTBmgcyN5wOcaNKG+G920BU+gPB2OiM7Uty4+/d7jzDwvN2JL3gb
+Axm6bzANysZ8iId+NggTpQRp6EXCpCC+AhM82eucHLtoZ0Ofkgl+78iHWLHVXfViFrzSOmAdrbi
PeuLp8n1z2ruiuTfFrsllQ5Owzsl0r3pANWzhz68fWbnOQWJMycPGMWxrIirbt75stNGRSxsJG0Y
m87W8Im5PgZo0GqvjC7Kz0ZA3/qzxc7R5aFRqBBizzQ/dPBe7QDltzwHt28MVG1R5W1dKQFfszyC
CO0qqkZHSE0odLtIDCjbvU7U4obKEhx3RZQiurGEXGUEVqUqmNtEqlgk5UIambLfRERhbX1os4lQ
8M8/tSDVzJCfIfSFiPjDY1eaQtO6IaB+z7f4EZpsn/nAMmwfJhU+MDLl21KAqOUYWnFqn51ZTy5e
bHUydZueXWs4/Vbq67xqe62QvqhvOcjK4OZ7aE8C//vLWcMhFPBjbZJNZGQP34ylyPfmn+TyDq18
QfZHEqPfe+yZEL9Kpgj59zWa/ADObLEPkHxrE+h3d5sThKjwBKd/3irN8jBVky6hgOyD6MHZrn0z
6hQMoeUGd3h5WxSLsWyr3QvIcf9HwZCEWgda8MTfbB4AKBpn2a8EA1qpjlQ/dQWwwIobg6sJ7kw+
B4tb0QZcskd9H15w0knFydWkFoQvMTWkmWlQ0PVQ4HK1razZykqMqySi1HKosMZ58hn2VBfkJ2Xk
sL/fFGiDL4n+ITXGXErOz06p+94sxjj8QgJIVKz0MtQhHw0DtcSG0v9mcrIT6one1coqTOwXnPRk
Tff5IY93x0AvMk7beZOCTE3TuhGXghenydPv9CMuddATK+CDUPM2773xoSEIJS4OEs+GFfcE6/bT
c+GRtVO3LC9lQ76Fwwvk4cWZv2dXvW37s3/bXzOKFSPTwmhBy4VBzDtgAKHwTgntPaijn/mabscz
4fOYb5BkkB2fLEr4X787A+oJ6nXR+Um1GLIVjapc/2UDMVmMmroR982RTSsk1YGAdYA8ZHa9auxj
9VyLMq/8L8f8XGwFEPZLyHu6REP/hpYiKPSagkTcqiQmRWpdVl4DBnErL+jgeYqacnjY80tzv4Bb
0x266wcL+3Y60omovTB4gyx0NwkVCDMz5hPuvyJLNIlIS5Hv+7xIOaR4de48nqz9zu9px2Dbu6/D
TeCgmzRb2sDPccLzBvjtboLvFzxdpW8enS5NmqV0OmwKHwC7JqagtYAKna84ILVbX5U6WOjVYjzU
KIfPxhXtJhitnoNct8lUKx84gPlSc8qA5SLTVjsaLwdRWvsnIBhH3tc7oABCssYvowS4qMQrFMTv
9m24dioVSfTNa6hmSkDACsMvoSXxZENAVHqsifTPkA2ryezbz8IdX7TfHlgvszhXI+QofUd4Vh53
wymvpjrC05R2Y9869VIjl2kzD9IHBsZDUKIjY+rN0P0aoX6xGySGiWF4+fSoXLELZOulmgHp1ijy
75gFArSiEGIydfk3dBMxW49EfzIABGBWepl9XDK8dDkOj3BKqpGEHSD+1y/lDC9wvRe7lGykkPE+
DZOVnEV2zN7hcgeISxaPKjfcpBNHhROF5vH5Do47imoaFM7IewhwgIZe0jIlIcGD31Y9VJHEXyCj
vOwDf+0JbQ7DD6Eu78BWxRP5/ae0jbZ4fIUEfo72HcbgwxcNHTy3stwJorPfZHYUi+/3PQsj2NqV
+gHExFCu/Hf4zBxFf7iwSkIgJhXIqYS4qj8YtyA0b/ba6vZWyRMU9/2fxFE+Vk2t84P5YGH+N8zT
TAgLVO+pQ6qvnG+obw3etZh0iab8nsi9il5ynVvMUes9fbWOd9CO+78uZYqabndRWx+84h62SNMF
1UPrUTKMFpljPCN4m+jU2HZOOl9PCUzp56LZAnjRzaVMqCDbkW4a7rvmOuE9hh+XY5VVnAxzGt+m
t8X6HBgOWyCj5btA754yiFfHiV4l2iJ4T22QBAgZxkO1NLJ+VahaGpDoCC0U4dxTLosXYF/seKsK
I6O/F8+8pN8s9te8lUBYr6lfpKw6HvG23wkuKTOaok5ugvGONSYd6evih5gCdjA1D+5Uz4BgU6Mk
3AwmKTWmnbgjPLZum3+LEL/Y0dnjScrEM+eZ+ymk63ED/7tCrZ9HJuib1euJuVx82GH3IVW3uyXm
BKEHqADJW2bsAqkJXd4CXMki7QNGaZWyNgdOF/AtBwdCfp9ZQqAxD5PQS3RbbSd4ngzftWDLnhEr
NRw7a4wTuSZC8O2DJiEVzf3itKXU65eWnUsTVAImV4+ps6Q+vIoNyie99HcWQovDn7e7Gr22cJnp
AQUfXxP+Oqyw2QM4jRn5NDIJr5C0c5lSZKjEuMA5X2kkRscbN7b8u3LhxXILfBxgJerr87OLDJeU
RyQMahLmI/8vCOgHHH7Yn6SCFxBEMX9+IfdMdZ4cKCeM3dbl268Ka0mQi04DvTVckT0JxJTzCwsP
wbc9U469L8SSyi1BaujBpmPimh6Vh41p7Ol2dftoiGg4bJ8TZIEzKL05ErrtD5CLbl5ysYjMkZpT
4zcWQ1VV/mgRWofr04exZUYBJjOaFoWJbavJwzUVEN5OGTfNGeMc4nVnwgR6rRa9KSMNV4403PkT
bnqwj4YbVmxeT7KgZ2x4u2pbl8hXiLUnTu5uY8y6pXb8udWdngDLYREQQHuqUdZzxRONmn3irLXi
sN9qWT7FrXL5vewxkCuklKAo++hLUx0/beED1AGQMJmIXlXapiJy0XjCz4sEUAIsZ96h9yjegL8A
MPjlBqZ+RWVTTxXjYf257zceLBVOsnHdtyNkjtkChGcgzLM2bVNmNUEvblOTgskHomipjO139rxG
yK8hpCSJDErf9LEGJMgVRXHmR88fYFfdWrcqufxfkZC/x54LcGS+JkhOOdW/tzkC+VFZ9XJIpnkI
rmShDmdQ9ZlobJB7y0DL65o31BBh7M91qf1LqDNp13AGvHthJ4yW+GIr/X3avF1w4Q432jM7FN4l
2Mucj3o2CQWky2HIfnN2M/U3YOV1gdWJwr9hsZw5LhrlIm3hWASz2EW1rKDjqRarqDVxBgMc3wwJ
fDzb7DHRyH0dqOgMooki/Zsl3fGEXpatIGwihNGXsTSFR6wTewc6I+XOQoakIhjTo+V6L9UGvitC
JEcZrAnNn75jKhsu9OfMWcgED5Egr5+yJWPQHSwh1BGPIsHdg7dmAVhRW+mhXDwPZJpp6txYESL5
HaFy0lldxnRZ1nUYcJ7kElj6CQyjoAWfCpn1tItZvJmulNuoVmfsDyS4sZ1UBuRKnZ4uERwWhgeI
5zFMUtJGSD8PYq/ia7slvq5LF17pcZymjdujDmEI7/55PnQzpvhDRYQki07gTJan7anSaZCZc8zm
70G3e+BnY5xZdbbpqr6DN4ivZDFur8qw8xxb+HfD7Su4gXzbUOSyPQ4GBZOqxCvUKeMo4d3qwhQf
2TRG9RD424cO2nl+ih516y0pjeOVy65zMhvbZhzcQoz1pmKGbE+AzKImdFiiobxwE6GZemz5Tr5C
qgudJvD5Byhrdbo0HeulkveLcAyztMVi6eAtAUupG9q8WBVohFFksqghKdWFQoy7V72ioQDLOmzY
EOiooIB386kmI/oojv1QKGPkw5g4y5Ol4w20Y9Cqu8b2iD+VDKdMLbH3iywusKf1BzZNq57DBsmd
C9AK1cmq9q3kt9kazWSaDuf9O/MukQBQmohxWwQIbTxYu5/vtox9r0hkG3xUcsGeQSmbwV/2gUIC
Utnx/6xxAXnu07VRiXT9eS5Nn0OIo0orwp6yNcyggIvVrV0UEbzf8m2yub8xIwNMUDFZSjuCSz53
GBXb+zfmfuvuZSS5blUyU/YKxCLvyEX35zLFZkdMk/F4ZBdMdXOhb7uBtImhdqQYDg5XmqQXiv/7
aE5sDR8DB7QjzF2kk4oEcTv71bRgDtrM1Vc06uUElDkZz7WvSDljiBn8TBVEReoQxYSwtRxlzpza
1QZuH/0tAKk73c8ITtKLoROApZUoInhX7gCew2DoR7G/rHqwyHeLpcaaHGgbFnKcGcpfKpP61XtO
EotxnlDGN50X+/WzmipEs0wm4l6j8Br9bYJ9C7tDHctq7z/Gu9Vy4vd7KPPxO4MxgRSTxPmFUdul
lbYvRecgOI9pptIXez9bWM5CbEVxBVZqeh6j3Q74U8+rXaSOuFcAskD8iCOKG8x1V9eMnTukOO9b
UESfrUTWf6qab+mvsx72dZW2C+W4LLE6ciQzJfBbtTkZJ6GCl7RO66Ee3fkFHi5znAhmfgNNccm8
/QAD9mJgK/CMrPIqUa8rNEMGgjqTAvXpRXUXHTf6w1O7B7TnT31ERLSrJ7RD9uzY8h9LaHccddl6
2CWB772ob/GySd/a5PrJFTgCWpgA1bVJ0d713Y7J/cGVwFDD0DKuqjDDUaMa9N+LrXJ3eHiNLBf9
ZcI+rg8pHpxL59dPDHi7AP178OetUvlIIao6FvSFcCGIF7eZ8svf34yY7p3vZjF31fTXefSuFWmX
yadFabvCIk5Ata/qko0rhu1oFyfUh490Un4Y5QmmTq72CzJa45onusv8QNWAsqEaNjoYWVIRIgDZ
0bT6Se6uXXHyeguzTMRu0QRJMJuZVXOXX9J+oRx/48i3spFvaxXX2x/EMVXqrne7VtcUuEwT3tcb
gf8LenwjA4qcC5RVCqHjfQ2GNBiSRfbvMXXNk3gpCfjwYmzbAHMuY4uLwl45iYyOOzV6vHQQdb4s
6wc6oEFoVv0w+WIU/tvAry3Xgjxho7QeFr1euxGc/6tlSwPTGRBZUVsLNf35NamYi8Xr+BvFQ9A0
HnqQkMSJ9IjdX18GYjyhTsFdgufpQ6slqoZHj+1rpqS7iDNnphhWNpoWbJbRdfLTsZe+yXE1+qqi
g6SftSfW8kH/QH3UDpkvp/Yn3CMKgMHttWM6keRu3k/rKyik9ArBzYU3RLBAHek9HqV8KCOBeHCq
hfQ+qDe3KH8Ju800ny8zAvRd2mm/NK+GJs1jhdH/616g02rytVrpvNcDdcX/NKLHpmwmZAzhRKz/
tqLef4nyBM2Idvl1ss44eCiVWdte6xNsVGiqUPbdAH6QKrJqYIv9Tvbgy9FIWOG1TBwXMqDMcaFl
u+sX2AKRpGQXihQSXo9T9r5OC0CsqtSWv2lFbzqZANLhqyc5OJ+7DAryf7euLMAkG29HR8LV3JRc
rEgMn87KSztjkH/27+nPY+qS4QQgHmLEBhOuWFvCMOYj6ULWWsAE2jZb25/NbVI8fqejHYXCiXky
bhb/X95wjMHHOakxGZ6I+peQJx1cms+WcAlmBT60iQF7xefe6V/52x6LYdllb9wq2tQAglkdSg9O
vMDzBgfXLe0XrCp5MmKRwhrw1E+yTbaN1tg0lgTGob5A0TkfVWgl0rs6ukTQ8OvEpYhDN5jLb4Yn
fLf0LewDhijvij04an6xDDdN1XCj3ABf5ZkxuYG9unsJPtVBH6Njt3YgLcZlb9LfMOPJLc4VAfib
XuWDemJLFg77bawEd/64ZceXNVGlbMY0wp6TYaiCraNMrB64aK5UcAvZqmBvIbRuuv32dHhTbrwR
K4qmjmw3/M1bwy1xUdx7skCbxoKaQjSy3e6f3mG/0A4HuTgCPafYHkP8mU5A5GOFT6Fj7cFid8Hv
4oqwgK1rtbhsr0hyJuSFKyk6izwvDKhvbZnuuVFmRNJewWvrCVbYbA5Aj6f+7mHoLLfoIFuTdzGB
fFImRuLwCftS3bZqrItXV55WhcSOJRlqWh/n3KkqcAccxYOKMyiN/vhN5Nr86aQnrWN0RNT7MHAj
Jj6r2bLLLYJRDC4aOVIS/hDuNA9IV6Dg2dN5JHd9BroJgXm3bXQAaKqRcy2cuBsptMY6qycw5ure
zB90q+NpU3drmYs905747cJwjdeolVk1VcHMBFI0o1plyd0i6ElvJPN8QSODVSl3W/x+NZEjPYWV
i4DlZfchhXeuSl1suYfiAWV7ECRJE8GzKOCOMXM2tSGHlDJc20oLwlihRSfPUbjIa5xjCFtycBzF
RT83r+eZeGwmK8A91NLtyIk+YPmA8+gRCQbj2Taovh73BW1zRRhslcrKUvIZbbiia9Q9H/HExBWR
s7Lxnq1U/AoOQKTz1I+dlybfqwN75GERf+BHeEKPkFXG9W/qXiwG/V8aPCo+75QE2x3Rpu0P8DIf
Nfof9JFAM8qtcdGqYMut3XlH0pJK0MgynV4sZwzBHO3zhsDV9no1b95YKrNVn5DIps1UqAfFKTux
qbPicubPfGhQsapDh7zd7JSMpizwHzvSzbuspRdqgfq4KmsP7b78FbM/z6ShXNDFPpu/nfjzEfDW
bf/XfJIZIRSyhTBiG/wXC68LOyYt+sceODLZRzeZ50MOCvGLdh0/WGoDUZe+iXGWPnx3sM+Lk2ue
pKg+DpDhSou5RdTUQT7jbIYddFlVFVYVHhSdSgqOANRhUbm6R5XFN1Q9ca7F6uqZJV73PbUrPB4t
XeWo+2TAxULqX386x2Crh6dirUdqqoLUQ54g8TggQOgLQGiVxNTudcDnDoHSjY1l4rxL5USNl/Q7
IAuhDuboqcp1sNL6DyGyghnJqkV4vIgbimHe4KAe1PqWb54xl4MV56Ozn6+sMx0Y9gNtnwX/lV2l
JrqP3AgCrIL6Gb7VHlCtuUCqhILM1VjvOLr4CaMCr7rcZmyTnzPuz02Ze+CPHupHWEfiZ+epxuxI
64OwnUWrXFhmqRplKrGKBjKv0vbTxY2C4R60AYC3Hp8gNlsOz6mT8FW0nusgB/rh9SWPNFdZzEe1
qxDQH0myI0avKbwChSlLFyeNSmR7PfjIOdyYhl8BP31Pulh/PHKxoK4ie+KMxMn9QGCnDNIGalVd
oFDa38+p4saGKT/ATF1AM7VvtRad1K3h5ZyKdQkMA4nYH5V/UKXmHvSVCGHDDcHTW9b0UHV5pyrq
EhUlloL0ezL2+n1hBf93cR8X6eyhg7sm8AatmLvg+7MPDljojqRdvI3/AkjCkDlChXAOgFyzRlKV
O1KD0Iau7x4+GeVOdpod5Qh6mE/2SvVqMralnQwpejMFb6gpHFe1CW+OFMVJ3mf0NbgO31XVGTw/
LKzJuA8ksuyBcPBIHHei+SDQwQw4ktEOVVrqkNvx5qdNWE4UJFH2IDM9fbg9Y9Rq2L0sI0XH7LPz
sZp6BWDqp3p1RBBJXsN7GpTvNtJh5VUhNL104SjprvhNPPirTcvjZoOe7joBNm4hCYjKJ5iaTepn
C/N6ykvncHgLpyVybU/fS168Enx+GSeVeDAcTlQoiTWUAMiSB0czt7GoibmRtkThLZ3YGOcyHh+e
aKkT3NPm1TMgBZDHRU8mi4HM9+sL35hEbfjl+zv0mqa8qb+LNxHQt6BHxhQbMlevApySC0g9jd0t
lsP1gJ9NrYs/L+Cw1oAH63Zv42cJDsfoDeySB7DRJZEaFaGTT0DTayRYvToL77FpJWb5Tyd2kvxC
iR29sFA1xgbelZuhKBBdCRAbeIcfarHrQMn+4764BdSTrIq1BjrpG9AvlZfKJGkwbovHFdjwqu1H
Zn2JohLsGiK7AHTZkB2fkbev6EVm+jAZGsPJJjWkimhRZ5LCCyrPwILXPSR1uJfiXQEAK8XCyIIq
ecnPmZqvFOwLg/1hJ5ZzA5tJXXAKETFBjwSYZPNeK0jmC96nraMk1/c07j4I5XzskvWHcIru7wbS
K4fLd9RFYi/fnJrt3J6xUCH3tUt4sDi3824DY6qmGPl2a5WiPN/GSgK6vmwoVR8WhEqUq8UhRqo/
h6X/vAi9YMvt2+b+5gqCClSRQHeABfspg1cM9+orejJQinoRzc/oHyiH9CU4Z13/k/0uD55/3oCE
a3qPu5UkdJOYUdKbEC3ZTTF8jYhqhtWMSgjrpcpCCKuJFeQJ1Z2KYw9I5HyDzUw2BN2E1p75C+L2
gShEZ7ds4alL+Qvwh8gSoTs/TxlXV4jq1WJbjQCumbEXr8qbu0Add0f3MlkML7MnwQdqGJEA9a23
tnPxDoOV39UoXIj5I0B7kDMN/KcypfX2x1Kfa3k27qYYZ0qeSD0O+7aF1a+zB1PPLa5VAiHOatUY
AnDByrIf5DCEaIDeYRog2YoQkcD4j4KVHHD8d6uF2WjPxnLJALfIoul3UL8bwUNi/jTErBTqsR56
b8FVJYDVk2Qr1gy5Cvm4ID9UeOkRvw/jV5swpp38Ha0jubKXF3gWN7fC0Uye2jU+PHnFAtCwpsRV
AHcJYCahHvn5l4dvDQXiz49J4odQ4rVB0jy8IvSKQLqzc7i2bVyKYEG+NUSdul6cDcFxemr6gccv
EBtJeSBqzKX+kxpKBveV/JANDWSA3WfzUgQ3aAgJIzrg0KVjiGFOAdPl6FMYGyrYpHg5V4LYJvF2
3af1VYv/+7Ts38Ghw2I5mIKbZ/IUoK0QDHcJ/VWSr35a4m+U2TgWl+Xn5hOvUd6DJ1hEiN0wPq5q
AaF8fn+xd7lavaiZD6MNUtWm4SkwRx6GQiENKlTnvM60uZgs0PKioihJIJbJGeztcqESDWT38bgF
PrL8LgqPVKQmsroJnZg664Y2RDBpM0wV4iu3m3K+ZeTh8C6G6q15jEjif+N/PDTYfhYrZV7Mem0j
aey/FvqDlB/0r04OW9nZ0SEWDWQlZO3akNzKueCYJyccnU5L4GZIimeXIOf8ReZ2TT+etMpE4ZVW
YPm9t8J9V+WQM/2Us3wsLoF7v04uGmMXwLP771bKHuHt9hMUPcKY9n6523hkd6g3GliBIgNApXMD
kAcVYy1Mlk1qVhA0JwUpJgxOAgV9u0DX9JDpwtqERLpHZGraL37c4UcksuoyAlJv9PSgkPpH5+r0
v31CSlTZodDkNwQUvfEIEnvE4RXLvpSiQTmD/RYdxQDKKhazqIzpRsn+nM5Za/ZkCh4hqU/BRNLM
dY+n1XUEtpuUU7KimjvTnbVRQYTjkZLaUvtTmBo639Jayzc3WcG3V6Wvwf0mu7vU496f/i7pM+PF
wDref7jANfHBSC7vuCf8g8ppxuKPTZRnhg8AXoVUHRFn65plk0VwCGHhXw7YkJ8nfCuVeJUqzsGt
+YEgYoB4ZpFL1is+4pJxoyQuByLlqoPdLgJmYASomke2bWKBD3IcVBtOuYYdXgEX36GDMsVVQvnd
exLSRt9rEuVNyadHeuJBhPOgH5K57nZzGb7O7QnMel80gq+viVB7M+7U5a4+C2fsSLQV0r4unM7n
UUOlru0h+p29vCZdPekAdGuOBleYCISEVxBeiW4Vo1DywA06x9eSkQb7xDjoqUT84BoAO6qdr9bj
IScLs6PHjTiUcQCG/ZbTqv0Tb0CwLn7+RXN4hXmqyBkMDjsQ0aGTihkD12CUhY9Jqwgf1qOgIxj4
LsKK2Xd5YoCkmSBGf5MZO+/NPU+TNADC3LTf4rwBOXMnZ8uNzuzp9U6dF7K7r742T8V5a9LhNYVy
h9KjNu3jfCZwoYGH8hVnS6kCs3+B4LpLGLihxAqS9P8YjYdn8mDFcQJFFJvCPANweoscNTwKFwmw
vn1iksLKgClSTSmYNYzkKOJ70cuS3kKeMsFD9c9WYy1s//MORobzGsuGeTmt2FbG273yxC+y4n0b
/Uq5d9PWh9Kae8ruyk92TamU+LBLGuL4cgBw4BTz7r2lKgtImWKj8pbKjXagvSmeKvPXdbRNDRLj
9O1QiT+h7wEBfygxuWsY8Fy3JbEAs4rKThNzfxqctYFBeN32lOhYu5m7wP048MuRry3W9nOjTJB5
EP7VjbMk1tYkP4xYfrniCNcLsdP1GMyo4xiG6f1AhMPIASgbxu1MQOeDnv/D8egkGTWPO8dDiJxe
FehCdLAXGW08Ja+WuCnA4xHvntreqChnWCq4dlSsbd+ROmDqrQGjxsl++5TyaTcxmUlu3ZW+yBOt
8XIrB3jQN5oV1pJTqGqgDxxUcga4IdwCrnEYPDCpNx1FukcCiMDLN2OzpRKfDPBzA+unJ3Cve+AB
z7J/NqKmYsbA7fXi9oODCBy3iMuM0792pQVeNMPxERcrvPD4oVBOROBRFFUPa96qLcXG7t8oGphW
ykjZrIUmagaK8YiOk1yBAFOGcgdUZHKWGuQbidnUn36weEC9/ecVzw6BEB3T87WGvTLyonwPUTs9
CSq+yB1K1nWm2ohIdp65mkgS5zKJJ4c7T5wNqUoEeCjUIIZcbo+e/iUZ5Wu7zfj5D+1ar0sj68Mf
GQ48rwjVdiorKWoo97ydqB2ydac2VU4JQ5+Q8Gs5jmU7yz50DWZpxPA6RbfSsWP8cjiy8JtXOjEg
SQ9bHm4x7loqgDOkdPPrVX+bJMOnZEVC8SvjEVZ1n0MSLSLer7RYYLxcnxdQLK3Fo2w2Je5Bhyh4
vkiPyVvHVUH+Co3DwNJ9vRO584a2QD9tRqoTWqtWji6Gv0pM8/HCVQFCgQnRloJAcEaYD2V/mP1V
hbIiyYZaWXbIPlS4Axgds1HKydHMGenNkgLQ7gM8MR7qlDwfo1DvPwLzrKLJCNrWD0TNE0ZZjnqv
8S0IhOcY7e/ln/2+Dyk5fKnWgwrpo7hiVk+gDIWApnZBIVWK+M+BA++FkK+Vx8LCJhFxgjxI2H6f
Z2sAGBFfbP91UC2wGpQMl5TaDqLkX42IVoHXpXgl9DFrMyVtxel4i3msnQYP+oQ6IByNXqh3Nbui
YU+O1WdOQuju0ej2+tfzMZQ/lnh/zV+dXD5KM0ngfm+NYb4/QICFvZSmsOZ/BBgbtyGNwTNGebHL
NiuKZlJaCv/0cvolvTkE2I+ItCte/gKwX70iRMcMJP2mQ7kGd3wgLJmhGwdwdoc4RXSpuNUa+2Qz
0ZciPIuB+FoNnOw2gsgCj+4HAbQx6/HsnH6i6ONU+dje2JoJGd5pHxgmdHpzNlofDXtcf0mkcdgy
Cc3RMKD6GHIZVFLFTXWzqF8VLprkO7sCdEYn/DNtqNOJZfLhAGWkaBTi+kus7JCas3qWzF+xYfzZ
CF5ynZza8h88smapbkLUF9pw6FDe2WTpnnS9jKjRiLG1H+bW4TVc+eNABxqQeiqRNTvV4/ZT1QF0
LwYBmxDrIjbh/oCXoPTG6pZ3IdgclvIRW0FGPA0lHX+zgvD/WqKfq+dG7JRcpDsbr3xt7r8t+rWp
Z/EnVn9XJ9vVh6WS++iYoQTFG6KO/94i00UvhlJwdX7Q+0kAsdaD0RaET/WP3FGeKf/PmLCoq5s5
CkVhUKen1EYRI/2se15vHNQXZI4ufj01X1nPyOm4u+XMNevRGQxHccMw1Z1NXiKba3cEDypzSzJY
yrmeiW1q7NpPP7evsPcbu0WLwz9JeZ+of9ktsiyeevhOMm3Oju2jza4YVPmtGy3svQ8D6TULBKsX
MwaTl8Jx1akE1M7/R4Nc1T+6bQyT+qwj1LMDkXnxMf8swruzi6HzlOTNedUMBc8oJVp2YKdIzo9h
DcjlzzJVp1n5HdpEDKaRxmcueHuP5IRKFy9P6Hys3qkVGrvO+AgSfIS2ZxJzvjfijvrGmU+oidFc
pg12eY0SD+AgkFc6QUUN8VQOlqbGSN5MGNW9C2P/Mr36gJA1x89NNs/Ku6wQjV7wo5SuuBC2nAYZ
SiaS4Eqbz3O05mXVfplRtVT0+AnKV2pI2uCP7CcdSbf8NS9c9ASXqAfmTCIuTOFr++KbBveSLjne
9ierkv+/em7MZvYT5MVPUnoCXsokqLUVRuHYYP9D/JmZ4OF4gVH0UpILscWj7BwBYmw6J/xZe/it
m71a7+rXyn+u6CqCOWrjAK3/TDJg7o4vIe37tRhsv9KolFFvSwAPp8nhtV1NcB687yfqE1yx+vhR
SWzBTAPwUZzvoM+dJ81VctIy5/nAsBgSkP7NwLlrNFFxZAloggc5pKYAWlQjYvij/HLkHn9d/26w
RnaO2CnEBNi7KXtjDRf+0A6oL8R/r0OEwscrAspEWIaMyQ4EU8WPfQLVeytHo0YIAvs4hjPIxlGf
IUUSp709Wzc2q8N+846NyAHdZjHE3/r/vwA6zrHnzcs4Bqr0QQoi/OxhmE0n1cAF9UHboUSNTrsi
ZzPFdYx08/DtC5K3KuyKyIzOa4MhizefHKOVTbWkdzjGk37IMoufe79B8Bm5L8LRgtzmJKrxIeKU
DN942keh4GLSeSkCyrpTLeWFno9Nzryn+o7olI+3mTa+GXGoIvi5d44VmSiXe6J/K1ClYoXtcY9r
gsjpxLaimkmmWC6O/P05xQyQ5aNig7qGoXEb7Kdsgzt8MPqrhXaKV3l8pQm9Bk3G+LV3LjtQyPXr
CbBxiifqaVru4LnTbMwNP6RFbnPBw/zSSB81im5f4ffB4wro0GZ6g2cmKscTVje63dLLlFp7S5t9
nrgKWpus5we+YpON0blr9s9dPs63yYDYWopQlpT35Ibe/1Y5mI9RdX5l6H/ytVJoSCwuniQMMobj
hPMmWfsNS2hiPOpNIKR0y7JDEopStuUiKRd9pQ2bMF0P2K8HCLYZuX8+j/hQFBteOe2EClohNSEM
VEQxldA/cQQTG/1OhLWKJHCwbrHISCDxFTU+nPb/S2Ao0VAw51Ln7u08UgaFqoX2HETZ4Oda98J8
eBSQgs8c6kyZk6++FUM5OAB3ftSzBsT7RandH67yMiAF9JkAY4F6H5k8F+J0bmJX7PBBYWrCsipp
3VBGCMu34KY7XGTvVOlQzqvfU/7yehdAb3LRAHkc0F7iH8SemNRBKx+k4sk4WTIFJLL9ESSqVnus
wkpOw0wxIomGhctRb7jdrWPvwVYjMuKIudk+ANEb0L6u27b1sZIuGRjj6fKwlthYtLYCjQVjUiEz
5rl235z6oD2QUUNc2mSUDchEWctaFicM3q1yN5EaBTduDDR238VXaToPiEL8VMFb8wJZYXPGau8d
TsiwTsejmvaTIen1x90rXAbwJkqOty4n5ds5WtW6FjXjV6dBy/p63/so6cWULF+LmLkSlcCj59kW
rNwSbYCrSq78QV5nuImjIz+rthENg6Jhp7+ksv1X1JPSfRjqbcOJ91eFZEilJHyNkx1Y19AppEE5
9VQjArzgiXPoh5MvUuxoNJkuI2slSNEP9SMOJuig4LfwMEl7/HBSEFmqKbjXtjnzalDwsMT4vy8G
QUNs66v5MHvm4viv+t0eiDhiiY05WCgT/WW2ZUUJtoZmGiv3xH6F96t3Mipca4NlMfw47vjV8qKu
CA3MJra6TN1qx2fDEKcmNulYCYDjW4HnUc8aDM7Sx0MVgpjZTBIzP/H4aaFIcw2WfrKpQnZvPl8p
79CuKSEuWYeyle7MOZefOSNqN+44KPbdsCiQ/N4Hhf1WuPnuVkhoB6FGQ0Ty90Mlde/7Tmxd1R5m
gzxNKOHGb/ojzL7MadwlH/1s+VcCDZZfbRS0VB+eW1VoTmGGGRfsn6b47aJIgMjal827CHHI38+b
HU2jbIpdxjg+xoRaVKBi6xFWWRP5wrYDwcmNG3167WXAs7//qTJXreAqZJP6QSPrsQVW1AMdEsN4
uJL5RdsZH0YKJk7lpfWZ5yTEt74D3sdh0zAWtnWmvGfzAG8XL4+gi4BOD9Huq8y75YrBKyUHYrv1
W801pCsOFxtP4xqT2zt9tljqy9mjrQJsiI0ixuLxBVGMs/0/KKC4H5H3e0JngCyOF7Aaa4ECrqkW
SAdcql5HUVE/MCS6iz704S8Mg/VX25Kfsfkxv+J+YLVy/vtu2k5JBK/9CskKju1vddtyNiU92xMG
SUWiv8qMIUBmkPumz6CTLHKVLBwPodqPEytF39CZPRBTcPOuCYEx3E9Fy7OBF0LpvPKLpqTBtTwi
huHuKREyxz1Ys1YHeZSNWVD/8m1BBrTkJVus9Cp4m+94BRUondcIMN5HwE6eOdBVODImIhCL8x/X
OlwLez7vG0FWlLsZccxGvfctcBR46cXQ70MmAAWI6uNTRvLE44uZaz2zoD/iRwoQ/hh2Ebd0ADQZ
lqoDF5JsST1TzEQHpyZbKEkhmyeeEuHq0Xe5r4pxXf88eDB3dA5Uifx9wGY268VbLqQgCtHajTUZ
37A5a38B8dPn6b+SnpVNzsvhPIyIJaCIbd6rGcHD2rJExyar/h8sxoDQdW91U8uq01OIAiwY9scx
WNjmlfaeWcpgA/HU856eJB3hiTkYZln6vBPkWlal6eGIkIeLHVBQd5FIwugczz6QL9Kf5r9Ew26t
JxeXssEjkx3CrzFBtrKIcoYjG8QL2DvNCe+/h5SbrtDaAWk9uoveXoIZA4Jfsom7cMJOyVPJSSgk
AENpE3H/9hq1hnfhQQLRRzdBPxRUQaBnOoPPn4PTrTcdOXLmpd3GKQRK4SKOVWkmB4UwlPubSISL
WdyDgNtAnwm5UB9Wefeb3qf0XeN3vxB00M18zWKbGAtPjWM+jx547pum9msP7RiKuEavKYHlpBLy
K4XUxGfkfjwLrHn3x1It2qBzdJcmHrDjo05e+x0GIoXOlygfVxAG+v7xJTT1WlZ4Wzoa/7afvm95
ayNuR/OQiZgLm8k642c+5j3brdqIkzVOVyU9V0P2KxLG7Gct5vm6AEVDaLsMvyQ/o402L09xTEXV
KZZzVmk/yTbUfao9+sSgDqB6IElJ+lOTxsWeLPbpjZt6n+osQuuxt2SBFTzN6/oDVos6yrb/6iXs
muGMxLxjVIqLjpcSPQzybGQ3jKzo1I9oqwTbR8TqvQXB7dq/+dMV+ZtWIYvJRvHdq826OYkGSFsN
XGZxnPgAYyuKkawbEI5bBGaiEdAD/rqzqczO2M+8r78CixBoHXh7gykuLc2//XuQgrevWMpNhY4G
xEZB+BIU4ZjcX0zlFgVMlTGwE9r3hPYUcIg/NAM8VOXtlcvHxo487dQ6m88EW8EzqhLOvUZdqjjD
/JD0V61K3NDYvnIUv214PSKJSYMKS+0zOGUxlStRO8kVY0mZd2vklKgv+roUZ3JdbOy8FLKCZ9OY
aPvyQ+B3uW+viEwq+QiHixcysRN1MsL9clXX0HvNgR/t1UhnjMmpZe8ygviJLxZh5KIj9LOF6r3r
Dwyf+WsduURmQwE3Cw33lrbk8csqjGJtaM3EjDDGdgzhqgYo6pA5Z6DqSiDJlKGtss23K3IIgCGB
OjNL6QDu2OoSquIBFpvwEmwWf52Le1lMBbWPN0V5nb+fP1tEuYiO/amoXNENPjrMGFygXdlgKZGe
DMqW/kr5KKrybmx1STxBCJRW4RzLa+qrEEaIclVKDilaL8JpLmoG5yq3Nqo4WBnbQbFp1lKsYFjB
UI65iP25Jkr6BZ3nbltkgy9O1EptlrHAuXBaRdEGuO0uJ+BvDDG94sT9DA26LP1UuGu4cSXvSvS4
oL02uIxmw9B3wGsDNgvqXNRwPXReIjG7vMxXmT+6kkLXXS9OxGC7dmd1dqCc0x3Szlirgze3VlGA
OMZN9N3yvxZEn5uUECDPFR4mj61xPKyzH9hV1dCwIdU8ewIyucooTWtx8C+T2bqB0uwG54B/YeDI
NaTq2X21rt4wY9m5Pe5JmFdkjtxqRDi4ev+Z4Ob4Pi/YZL8Fn5daM4GR1rp7DtUrz6s4VBv/fFHq
rNCOqCMRPxkNMTvN4Eukf0bHFzvlZ0VvsuxGo9rtPBVl6kKaQZZlIf20QnJhCyITg2IxkV89UusT
haUQo/nT3PRUkpuhHVNKHQljEyKkOoci9DHQi+6Y4aYui1lF3A+nNSvJgx8JvnTcRtQfVTvJRgvY
056RE9OmpZjxaYlUZT7yvD5785qUuULaqWSUZWHk2BRlpFm1peYO0f1vpgj9UOTaIOK++/o6feCs
gtrvyM9tVlsaosi6VW4Szvhpebk2huwGUBcdKBsKLST5ScqhPZRQ48HunoDYg5efM6OchfP1b2ft
Hq2VWtb1/1EdNZ1VArvYzSF8kKrCXbA9qM0T+w/OTP9p5/sTqkTACxPErYdpB7flA+fQ0Y0X1mK+
b2rmsxppxi9XtWe4oG3cWysIwtqGcxDQn+W1uFLFQnOvrR3cj2lUA86NRrnFCkE3l/5vUY8r0bqH
bEQ4RtE/ho5AmfBH6nNLooiICAOJ16CK0sJbHXZFefsE/5ZSWifZJdaG15gdb9eHsHHrB9biDASv
N14iDWcALYVOHqxLqFS0ps2/+CqhrTqPk+RH7wKPFvyq7AA9WyB1/hwUeTqXGYYKcg77WtuIFNlR
6EqtFgFP4tIEyP7F017bOmA9PqAVE5CfMrA5+GYDU6mHbhaCDSI1C+qb36MtqkpmFto/mI3/raff
hllZja2ZgKZ3geYdZxDCKpScGq5usm8b6/3PDCnyFlIdTW3dfnFFjQQEcJs7nGgGJlvUYv2lmoYW
1kfmrdrGEvhPDGGAjfoMp8ezYnIsOHtlEPOlZCyisPwgWMlWmhRdV2rnKt/aC9vABeAQmFzstLIK
mXBleRXDG05YNUiUxJ/5Z0c8BcGKfVPLLLgmf1HpZuWJ+zas0EPo9QYZAYWiwJe8AQl1m9gnWPIM
cqNOxeX8kOxvhout+YPhJCCb5bCgRU4S55P5JrlYMSOGiutei5btBy/4niB8lHrTZ8siECXvcr1R
VPjyNOQh54UxE1o9eoHSBt7rxJIzyTgxSzw7FfrPU6ELgSK/QsX9I4CGCmcZQIAt0qmv8MH7oP1S
SMAqBSsrWKjf/YKEQ/lbaa0O2jjoO0xGB1Zfi6KhfMChBvwQ6s0I0byRW8f9HqUz+9t94o+9sq1J
mteweDJUSal738UtGXuAbpG0CshgUaXxvEp3rxmg7gF8N5XhDb5pD4RJqlaKngsF4LzySCMra4pp
xAnJ6yBJbynTzLU2bQzZnPGTZ8AcwTyHtRb08vQtBxIQ9BITiL+ZpeN4zeEldN6kMwOUAOsSyIxI
h8KWuW2V0fg63CEb0JKa5+4MeL6cNgAzRZjYCzZz5AjFsvqhfWuUXmuM0tORqRnDlO6Cv1vX9lCD
WPnYmYJdFANr4QTvw85cUvNm1Uub1tR2flA2E/4G3HnWnqlw5gTtW6TGKRmZo4R/KIK/Z8OHasVv
ecCBnRvfeJlm5CoL76hTwt7KzLUkdPpSkga6zEnfcWB/jDFWxiQV+jLzSk+QN4xXDTpLkaWU1vNa
wQWzzpaoURiZoHGVbrQOzWsd5V1ZxjtuxNrZmKJ5YQayyGlcoibswA4N0uIuEKQ8WTrfVau00g5w
AKIXhILAgOVp3xYA3+EhaNTktn5rcY9K+dwemm3J6MjjOc4iBEfa2RUXKc0rUIuIFuchV545zjcw
Tej6IXVL+QFy5z61JcRyfwyhqRyMeH4vUu9L76jxsPy3rsQHay5Fr8N3pxebanN05Q8IB0bCn3Ej
d60PyUuRldivMdOa8+Z1otRqYIjKwvhhtHxolJd7h9+JlUucAsmmBq0ouLYj9YX1u7FTzzYPiqwt
0Kag4jNGxVgss5b7AbA8xy8OXSnStcpWN7AY+IU6YaaN7DK7nXQa8RiSzzTOVyebP8QG0aXJ/d/u
Pw2+7T+arnxXNqTR0fOExpIVWj5c3+GmHPPEds+InQFuHCF+l1hiDOIAphw+h5wOA1x5C30HSkM0
LgHv1JOX53YW3wHA/KGedNlpRxn7ihSffQFp66+45BSnPR8PXsJLJ4gGmtYuhqx3E1j5BNdwkhbD
nkc0DjkJ9vBkViJ8BAG0bt3y/jLTsNIUhKCYlO3dweeBkg+138CUySN3H0lP4x564OZgK4pbfXIi
4Pu62Gapvnz4nirVkdRHwVuu8O9Lm57qfKzwxmvkb5a5R77nYLb6NEPUbepOxo4pjdhnAJTtwEUU
41/Abm9d+UhecouIi/D1EQlA79Qx9ZajnV48v5sP4TUezVF9njXpnaqTQ+Iq5vNgz17dVBEpRriO
H/zrdPdxTQFzc1Qd6OoJH6kl43mgMGctqdtNOWneBxqGb7/fBcbBsZpGCKwue9d6BYvpPcKDuCcq
Yfbztvv50NZVt1eZ+eFsF+M0ec6yEIwowws7fvDpqH3GfEOp8xt3OO8pchnpnaXUmVm8sS9p5oRh
tCQpjBXrbR2pVzTrfZLLuRE5VMu/rtOLFfLavtAxWwcvaBSt7qovXGEIB31HvNEsGBhA1WzMsD8g
4apXr/cZqq11dpY+5V4S4Hc+BMiQa+5L85DfX5aoRxtuD8dK3YOqN2nVQUXguQs8AFOIMipbiXbE
pqB5SfeCcHn6EK7GAbscd1qp4tY0lskL3+JcCnyTdRu+Hxn0TzpAciAe9B00ghdqHyKbLOhJJrTc
QZS1Ifpm7ssKxmDLByeHgVVbLNiQV2PpY8qjkHdkn9Kktr5uoPcTKWoB+9aRBTe1NN5HQgLOlFvU
Wfr48k237LfvXW492gIPub6bvJP8QyqX89YXPWg3WOA7+qjpWl6JCU7fQ6Nzsj5KL6CGR9UXcgAB
WDy7s7UF85r3K25WnbzyyGAyDevTF20IoLxZb8rt0J3YUEEVvB8uq0fn9QS2VDvRrcTzOB02wbRe
gdYQCID5DHYx35/83IPBAMmSod10HEvUR4BTkBzdTC/W7MNxAOFDmxfmuRK31EHzMANyZiGBrPQO
JfNlOKqXuo32y00+2rgERjrBpTenR3M4TmY6Vbq7AMpFsPynsAAgHhztWt0NvDdPb0qOK4AMPjPa
EQSX3aDkztRhMEgrQIZAWqxt/kwhhmsMNYk0Pu6/jZ3SM1KQj7vsz88YzdT10VGfUj3V/fCP1qna
yJLsp92o+lNmFPz9K+vMjAo16zff8d6wzw63ukzJzzVgYwgGGmZI/PchsqvLtHQNVjOwidT2Imnq
aIOXdF8XEXAOcZfmG+0jL8X77eZVSzvCPVg5610ePmgt5gGBjNLY4os7rCyjtzfFmuawM0DpybEt
Onenv9hSGQV0yGNLtAvoEuigZIC5TvC0z/amLntnj3nA1f8UuDqDQ92f45s0i7TJ4oSBeWKI5GFF
En0WbCF1m03cL5XOzt8GdEnX/NgmOKUTD0CryW/h9RrOuE4OKja0/TBEV8egrX1NcVp6+GDNavnB
Q+Mlu87wcI8iU6XizIBaSXfXhehF1WE6+YKuAo6m8nvSfVFlm6A0QQxQ+IEr/PD6RjPTVsNX80Gb
aQT/nECRB7yrwo2jRHFrhVidHmDIlSNQjNgi1nXnP0nXsMFs/sHsxrl6ZuPcg4u1NME8UE+qCnjy
L0tzSvlG8Z93NkXuwgnm+0VS5EKfrlPi3qxf/ZlqULAEJU9v67dRNf5u8Q/RDHqwD3EfrjsuBfQP
AvOqNZGCdPxLo/jJunxKOyLAWlgDvI/XpeIYzwAy7RgAGR2KTumIPaHwqgR+5qhulX7lW1ABzyo4
KWSqx5Es55EfRIqhu+ULGP3x9DK0Uj/aUG1aTC8dp1dt6HzgCtcDGdtulrARurpfcpjaDR6iMSMj
+84JpaqF3RcOXCOIneF5JLTWLFzwSC9f2WqMYpr88ucWx+Cq5RbOpanbNu+ZyZ1dCAsjKtuhZ3e1
2tsMpZq7V2gGR8f8Wq1xttq8TgHaJTCqM0S0K7n2b8Gw43yXJuuVw8dAV+ZvQN9ypTuZSBL7Rdbh
lhDz/Wip6CvhmrmT8VZayJd1Z2PVL1BDafFhLWPjbyIfQ0YLUWv+yTA8aPg7nMDwNRxFuvrWSe6F
ftX+vBznfTElWTPx/l8qJEgWHLTuTHKp7ClwEm9biUAeC8nWdfHkgXkoOzcu0YU696XLODwFeCeu
ppxSPDQVoU6QamqHve7pvinI1lu8497wL0QzjsruBUMXOWqiFcgIfyC3Kxw/93SSlS97r9epmyaV
JLaCeOuCdXDuMusKs/VTY9eIKGoNfTLhocxKqmlYVtdBYL7jw3WubhF0X+jh/44gXqOR64W6tLxF
grSGDtWMGQqb4Wj7JE440D3m2uFe3Z97xTvm2AHrK/iiFaIyYPx/Ejb9ymDP2YFFpNy56D+b0baF
mFl4biPYtKyO9wm0OczqvyLrMShjIWYlhwqxAmeS1dGcbBVNraeTl/CtIGB4wOAnBB9TP/IZL/X1
ctBruZ/bQksJarSYaAxEgCIkbBVhevDy/gR/84OQFPKr2R7PFocjhG1ho++UNdmSvkwUuNNQKPvi
9r/OPD+1VLaSUsv4pN7VY5JxYP54XDrOUZo1wC5IjvZvX+jtYcWaE7yfLkkvMXIq7Ws2GbZMFLE5
4pumTidQjcH+qzfCQgi9Dyp8QaMVnDvBfKVx+yIruVsYs6L0+3+/MwdjA2PgId28hkJxdGCCU2Hr
CxaCJebCh3FBT/7/4LXNtwVS8lfiMGhRr2E7q2zM0aMo81o/NrpMjPBnoAdYJxwAEDSUP6RWXopL
/kZGTAG3vgIyRE4agVp7jta0vbD2wibE1oHEDiWmBrtOwu9zayZkUT9Yc9hUlE8j0WOnEdrnD6v+
jaSYT/WBselE+q2YLoh7yjEAYPaoR+xRqEhGXp3+mFIono1t4vYvxqduTZ2q+9KOtTHw6FTt7Llf
Zgu7KuWsHd9uS601exijXIZtjtuM06gK5ovHsnFnzUeAyGgvc9MN1iRpO2VGKlX4HBqRAQ7zMI61
UKl1SaFdpNX32j4B6FoR2QGNEipquZaxf4itNtG5igHDOiORKO7oHOAdNWVzaADFVkrF5cTFL98H
s8/aHhi5t21ak+wIwqa5BD2fWGcRO8gtTJemIDEKE7J9z1p6qnguLPBrlHybH9xtZngZUXiNMaGd
5aAY/QxmEwGeSGLQZeII6ZFsU108HUVJcGGbUgT/8yKMH2mIk/WoEaqw/IB5SjLDprpUbjzlmPCl
rx681PYoNNwxzALoiJqCkOSj1rBoa6SZeJwmX8cj2FTM+MqpqlOI39weFlvNykaSOdx16LqezBVn
I3UhAPp/vpCO9bMpyxaeDN2skoy/CYegU/uSdQiwmo5+LYhhP1pZN2jxmrXUT7GHe4Zzm7JaTnYF
zrYSvj3vRtNiGsOc3Kh8j/s7OY6bwWFVSnHf/eV5ZT6Ir951zBCcl3OzI+b4epUcycEh7Nzx4Prc
WWyY9cOZOwuHMmiPseBu8Zj1MfosuTU0aIN+hN2W+bzvRQdCBXLGZsA59WpXND7tmI4uSDRu1ywz
+UT05/0MMQQ0D5hE7wxgilFujblxNpUEbcmhf3ImP9zemAE4ewZ/P/EvTZhW3zKaDqL7xA6fLequ
oz5k2ka3bUe5TDpTr2ZKG0FRf5634kCPR9Hf1WIoR/9XxB/84R0vy9F90pfhEuY3jsKbAwuWpwdw
VxXJ1guEEQ3iNa7haY9xwXGRJDIqFQcd9pfy8+wds8hB0jIs23R5mTqym+14outxcx/vamG5Lwm2
vmRVk6xHEK3bcFC0tpwtJMi1MFTFP6wo9EOXz2IAHNw5PnDj2CVHqCYZzJa26urrEMtKSWDENYGE
ec4oOkipvlnP501MIqL9v70MRem0ZecaRzeiVM1VmMgi4aG0kOHH/GZMnDlAmlZvse2JYOIsLyJq
8M3ilPqrWX/nQ6bkRt2FCB2bnpjZg1CazCj7Acf8Fk36waAaoCsTgwoCb8+EQpqqcCYJvRNeRvpw
yoKsLZ4RalA6iUN0vmGBpK7jUc8YEiNkhyKUoLwsszOjuNCTKR+73vVCzNQPlAsCwsalkXI1Qspl
0NGRQZ/00rjGRUdhPkaqVXBVSJznjPZfR73oB3Xj+Jt5uJuD+VYejx2iAiiZ8troBBLDkNLzuGpD
FWnGOCVH3KBeyCNTU6EEcb28wTahLZr6VgTbpygXkz662WWya+5slD+y7U2JadVS+JPYS0NAyFdh
TbemSxOrIe27M6zZh/iBALX4fbjjTdkpx0pqBZUlNqb9MLqJzE5tkRQJpbf7kVov9Mmbvrfl8Rc1
eDdh5fmnBR2dlPF8NcYNU5OeM5GKug7dp7ks/Ufx26TLds62JuMuzEUoZYxSq7LYSJfQEY3M89yv
LRU2Ec2DUgP4wSg3blJp4mdyrTcw1W6MqMAyjlyflTpqYInqYYszJmIKTSJMVrPAwlNDlmN6ypSH
dxQvQlSyiiAoKLuzw/Znx+OhjL+6W4ByjUJ9sFsIcPHjFiVIxbR6n4gepO9yCR4fDJEaAdN5uPJ5
kXi7TCY9nYgUnpSMc5Wdl8/4SDgtDn9xqa8AVaJNpCl8dJXmSVRUjZXso8SDuFoZHXXFFeKfO/B+
QfWHwechgv5DAwpHdTR1az5dC1zFTbDsb6SxbGvOC4Z2t2r3cpZccR/8XjT2B5Z/CcjzX53Tb6L0
+qq+Wvhb0uvJlJAxjLH3kSmfSRZpPLpzFtTZP18kGxp5hHYXnhDMddAer//1DlAYdHEaPK1liwP9
UVQiOhdtPFWbUmdFdNKcmr1rIhD9HmW1E8yd0/LFjSc9tQG0rGCZqUvFlfGbr7vyJ/98uJXfoPlQ
LtxC5BLo2a0ioVlyxYZLCXCTVG7TkfbrKkSC7AfwBzcO6TNUFnEkwZYWLvoim8Q130tggED5w1SJ
6aUfLFhlPP0i3KMrvYecq9cTWKAPnoVlberZegztBHwTNgW690sCte9R2PrURv7CPnf4UluhttB9
8wjxn2h8UvHAvjYsFQ4tgMdBr/lHKAdjSPrizqj2A6MKGuUfu8EfOUwBY6WNpxSX9Ps+ryiR3lYZ
dRRMS630ZyLakX3WPxrBpk5LfXT3TWo4Z7WczvQbRhygZDCTcqSwkZPfkATb144rLcGcMilxrnNv
dXCbDd0GwmJRlh2LtgAbt5cluCreC744wpodYVUGUX8FVa6asdjGsf6zt+2bYc6xioLrVFWYdoKU
BRGPvfmE6MyBmdwG6hO3rew4Iv7qk/cmCPM30R0OmWPkAV5AL3aJ/WrFmd/ubqp/8yMiZ/Agroql
JcfcnHVEcZa4Hr9iOalApIKYChgyCIEWghD3pQfsox06lv0DA4jZ79v3ePqIZGOgSe6vi0Zqg44t
w9IutgVGMTjpTfndMN6acLf8WlY0jnUZI5F50/3njVPEOd3ab2ZMdbK/NTk0Ok7Rv6XSByU5uDKT
s36HwfPQpNDoV48TCAKMv+6PRToZ7Q6DJAhwAVXKYNbHcBS4sC6a5vO8nFLouWn7ffHeauLAJSyi
O8ZRRVd88kUfzFkHgZ0a23ewDCWfFXcJ+ARTdmC7L8NgFol5c8D91O038qPK0Ml/AR+5FHP2wW88
nzNKYmr19JIvMRhjltMYMHK1Zxd/Ckh+IrMypsTNonMLkK8a7Ncc53sELpgwDR5MnsT6A8/4hukc
MDZk2JwkoKoAZI2ZIidhzANcG524YDQ7UKSpiKsK4KWYz3fI8vZ/G5Nhh1w9aufAsV61UZWnrQfa
9foTFjHj+oJ2VyEIqSo1npFYgcD4eI5eHetiMYJO4EiBjovZ08ZQsVY9Q4bLxeHJBm0whQsLFaab
fNcg5ma+qtm/678KYtkNIUSLJO9h/bIg/Tq3bIS2pxH7EFzR+QnN5z/kKE8lTPNV4uOxZpHY4iwy
G8EKj5OqK3LYhkGBZuq86nx4a5fc2NQwONiH6ktpRIru90BWXK+Ivzk/kJwkY8607qQTdWD/SZhs
K0Z55IPoKAy0FyjW1uNYsszpZbZNWZJI2h70POiSxN64zJNfuNhvnfKYRwJ6MCWMUAMyU9oigBvO
5zORvRHuremmWpd7Dpczh/t3KQktRRUR+T5j1ZCqOvhzBD3IGS1gC8y4hvERp00MgtJfg8voysIw
DlCh5+33Z6vVWXoz02hF2str7bQZh4+MR0P3dGQufyQg6tSbqORxelewN4EGbXt0YcvUJPva0ww1
kTyz4YKHbL62FcQ6G8MJgXNVZIytxBfFuswkmldgO0q6ompl9B+QUnhhTAIuN+Y7se/8gtMLNMWQ
KEwHmRCCzr82Mjym+uyVhGKU19GjO7h2+UUXNYMnB2LkgkGMteOlogLCH3kLuOgdXzHmy1nGrZ/6
/KrK+Rpw7+TazlNgYnSeFbY+ix07teS33cl69NBLGms0huwYB/FpoVtjeXNDV1Z/KWp2ew6/1xcn
WJwNBKAyNmPhqxU1DfnJBdRLvhHWFizDsDXcr50DFqfU/6QGJJY+eR9dUWiHHYjBpFHMrzrizoFV
4jb8OTMgwzp6oM3Yaw/qsQIWBM3NVDDUW1Iai5MC/uowcMRbfU/hr2adfyDpQEC4qeQaGeECsmn5
bcOyOssTMqGHcqxgYiFMcx0bgN9CVNc0WvMW1jQ9CKXTVAFDgaALglYAcfcIQ0H5NRscDz4x8K3q
YrRJsoSj+GOcnIxfsyqCIfzUQ5RJ2uVSkwbqMhbhF1XpDKw0PiItcHeGELABCSC6NvbCXd7mB6Dq
lYJcs2L1Fhl9vIEc6p0QFC+U4Z4VtF4RD187BVCqTlOHHzCbQ4tc91Q9ZqpXmVYuDi3tfRsgKY1U
m6dEfExmz1cFJu9XDyVXHwWJFmfxr58MXyvCDvYFaQb0qXxGmKiRJ4QlUSVSKXwZgv0ZjQRicN5r
jg/3ZXHRD8rzr9KDbOAyEax1YA+SFHZXtlJn2u6FEc05sg+RRTm3//ge3ZxaNQctBtqVqV14Yy+E
2nwoJ5WXh36+76zY5wzanR2d1rgilomqs2AVShDiBA5GVjloUFoTEm/xUD1vNat7DFLOKutWCuBW
/gZsS7J/V3EWvueLElIhGjTVyjoaQtSDY59Yt7Zks0yFoBPn+jLIbWhaIqOT0yQOyCuQ0Nme+dEX
ua+saF1e+XyU5EVy3DB60XhULru4M4iExhosAdIR5P3+tdNABpSXTV5gPGD4iMvhSXcuFZKcvc6M
DgOzDN0zFy/LzZAedOP8f52rvAJVweqWHgjpqHx/Ury4DYZAEU0Sfb7LqyFf0ec69laEICwZbl1A
AfPzTaQDsQRXPwHi6adDKSIZYwBncMFW7arhjwSiFrjeZGZg/OjGiD0CWCeTo4QiS0YW8/9TfTEV
udbvtlWaW0WpmAraCIjWpfKcGLlLaTtorsZ4ID/8JEtvJyf9PuV4ilwaDqBs34mqcJici9pnZqn1
jxdvonOensHimq1+iZmxC49wSGM4iTVHjdBY5k0P4c1DoDA9miKCIqD+AXMUYpoiE1OoH4E0WidG
W03Czx3CtXJeMXmjEYM/Sj020bMxUCIDCeS5B7BwS5ZkQFpPPaaYMIFhmotMY0cjncf9SR1AvnVl
zG8TG1t8lqDDKC/qJe9JUzFdyQ73hEk0W//3hpcY01zwihIVavICEwnElT/qr6L72cB9FfcYngii
pNZUiFYi1FuPSnMLMlDpiesT/eX9YkOHWUBdZ78/kxwN1Zn1z1TKoTPxZvZgGb9Iph2cTH37a002
Fc57+BQYsdOa6Oxm9c+DUuBD3Io9ILDsQuyfFkVmvwKfiri+5bzy7Y6J/TTCbXNM3gzjw8E0EWFa
tIhgS80yb8B0Op5F6ByHiW1Sh9jD7rfaRgN+eRPmw/yjNL4r5hgMUoLEuuA6p4syv4+yL+YLmuQE
i3vLkCKGlSPiljgWCeH4P6aaFGByZchdYeZ9d0yuEujU/ObxQT4dgIXdW7X3eM/pmbNoAuetKAmw
o0qZHdR4TX5SuwQWyXzbywcAfidFCveYcwcm2/+4LF/1rdoH8E6kqeYQ/yJm67VectRo1f611iIQ
P8b5XKyPRnZVSU8lEuEt3mrrWb4077DTmFwW13LJhIdkoBps6SfL1TWcsC+YChz7ZgOlyaOfNzLE
O3h/Yf0tcNm7Yf+xAjV4xTrMqPvE3aXo1Gc01PGUhqBxVCxdAy0F5WNaheV5/a7JgNk9okFRTqgU
D0hofhUCLsGmWwjNYCjEC+YbN8dsq7+SSfBkGqEzWzV0f+HeZolvcH3UuotofUFazo6IUlLU3XIl
12vKBRZqkERiwr8wIRh5dE+4tGP3x+M1Ytv4j3iXBvyzYdEEcEat1cJlvydMJVku00H0gRJY0LSE
8CD0GWIqQsnyFZvYQkm0yu6R5YMZEhth9Hk3huY+hgO4PVlcpZICAo49e68MzuBZdlgL3zpFm+5K
GCRZXQUAXLSl8qgR+0tnyM6C8jLWKLK5XdBEUgF18OfXdTZYRvNL3yujdbEHchT3Kw9AquMufahv
eKJRl7sJGCkKDrst7iuVy5eCF8mFSG7s5FKqeYXOrUv9peLGMLzq1vvrUJOyPM7xMAa8f1RS31fr
bf6TFPsDU/5tEegG/aaW/F90EZsKUm6KIp6LBA0V1BGvd5tmhCHrbzewOKeT/MnheEYEgoU69I6r
6eepqm4MUE7hc8a0YJZAcA9kbIb80PBcDXe8KrLibY6qTlpz2ETTI1s9sxtR/3H+K97gAs6XybXM
9iQRdQNveXigtpBRsAJ/yTpJ3OmPnejzvSX8zRw4l9KEZ/jdu44rFXqryhNFGf5t2XljaBBgDwvq
ro5B9AuF+VQw6phEmGhW7myiYvutvv5CRkN+8VY58BTyreP2PpMB/np9ezD3uQ77BQRQsyyrbss/
pcgHAKwLH8bj+wtOdStpRz3yrI95TZjLbQ4mpdBdfSusV3BQnZ/urzN94EGgZMlBzRWaTCHzVqyp
05JuSNCxQ5hNnaZ78CbpVB3MiZcUkTGgTuFZkUYFsM3JxFNusEVoIToEULghZacGKcFyzADwBE6f
btU3bK9Mp0OOql+83NFuhbPrzM/rFHqUCTHYafKSqAU3Q3izagoqZY08afGvyd2Bxtzwzzn27jsD
8ymrqxPgcOE9HLOkV6AOBjKvNpMAUP60voinXiMgy0x8fsW5W0GPy4a6ml6sXMSp0EO9uol7BGzR
F9UbWsNFMRnaZQ7sYo40U8kLQ02Idtj6GGIDwmUvbpYyh9mnq/ni3DN/OqMMbguH9RN6Gmn9dWra
r4v36B303q2NjuvKKAGlX53jlyPw9CA33xpi9XyJsKV7dUZG5VeUj09CXWP11HwTZRiB2O2yLTPb
6n7CU9vdMKE04QGo8NEiUCwQNjNTgdnpXpCNWK4zyqrYageP1ST5y6nNr5EXiqAKjj1BnjGX/X6k
pj/g+CQWQG/BEvpgWV2vk+w3mRxYRG4H2dACMtS3Q1bt23+8wqNqSmL8d3/HjHa1uTJEDL5ia4Fp
705By9awBlxt0fF/lpbGBrS/YQUmrXhG81m9bWtugF+GdYUR9/N03VN4UyctRaBUY5FZsSt2kUPn
I0AVoJN59ZT6CKqTDLw4lcD8w+l3H+rVknyDI1sfp1MEel2tViURX9Jg2eFKkklVwJl0W0T10wzy
c4zEGf99ANMQHqnUJrmfwu2AEW0axXW2+GVRSYW1TeBBCFdti4nhx6tYl/WFV8Apyya42P0B9X8r
Fp+UX4EWJihxGk8c8xDTiu3DU0FuhSMvm460iH7PWUVIuZGgIayXaoOB/Rn3xyR388TF+ySo7Ezg
Yllia9qZy24XYgZ1UoC58Sh5IM+QfYPNnehrEo06CVw6GzIiVoKTOMfHPis2Sw0ouaWJ7pJPDu5L
5SiNcbEERQ6omu2rqYpJxUAOb3O3ulJH5+5hXphqG0et0VClRbX0kD/VVqf4sjVnmP9IzVp0jAjp
W8zZVYzyWkhbO5l9n52XQHPi3tm9nTj6SmHW1t5ZF+cRcmSzktvsLGxMWH/3UkgENmmiA6j+JTAI
p/KbRqyGDbCyCABevwSgs70+19UEOqzYG9rosRDDhD65YgI8puZwgpzosTt/rWe+STRqHURYS4B0
bGIWixLUaBZRa4u2lpuZnc2addsmxjYH2gOLl6mSuEvxCaWUwkGdIL1Mt+bqsTSCp/WZG2l1iUNs
m6lHcWHRMYQxSScCYP7wlD3QyUyMh2MjOOxcISHNBcHkNRSp8633AY0kr/schaFNwGAAtsoKJfJK
Oqqk+ZZmJW1diIlJokRLmczTeo6I4h47O3iuZi/OeOwVtUfcP4ch+P9uZaYHKTe0biJb/QjAjMNG
38mO8xbAYMW4t7IvmYXd3ciDQ233/RPjsL9M9DVshGlm1tfrEpxYycQSkWQxyZnhVW+PDMdJCp5L
XGRawQBM64tqKuIC+Okt+zflN8mcTvCrY+Eby5vtaYE5bqDrnI89oqV5FdLjZbk5swcfU71SHLdx
+rJEEn0DciaTB9obzbu4IcJHDVSlm7xus5YV6OkOvNkR/JLpH4k3Pc9jyOenhrUgLE3KGUq+fojb
nhX+X0FhaGi9CxLIlWx54wJNVVfU2tG3kDtzLgVQ/4uy3y5dZk0h/pFO4lDiGZbXKgFjJr7zpPrt
j3sUPabumd2TnDbibKxDFCXGo6BkfYEKHkhAi2iut3nc7WoF3jnT5S2o1zTipiAN7Q20rYNRY6RD
3Pk1NVq8i3BEBrkNuq0BZQsdbq7UYZtZS5aBDhWE5ZFVzVtUxAhR0oAsRIuLqTmzao/6kIdXsVIv
/FiZlOEmMTjsgkPMZPuXklB6mHUv6m12UWV4XYLnvgwFRSvWgcsW4I5qCnb6yqFQnRJWJwp+Joz2
t0zn1KMB6WRhk8Ub3EZIi0Scx/4eiPUQtCFNwUBmiSQvnYGH9WzgvscRTM76pQBeJmnaOY+tOUTM
7aCfg4Zr/Zo7OP0SvQC0nNkV2GRzFVq/IBvheS6K4ZF8Dd48z/A4vx2qc87onxgVF27NE/aLIlus
ryH/jtSqQ4EdO7P1tvcos6d9ciAUvoIoCzgDzBJGTVycxLDevcglud6WR1mKIT8r91g29bx/Ww7B
/hPxqOGRqow6susD0DJ9++iev+PjJ462CeE5Gbny6a/WrO/4WVJFBz3ZXbeamboRRUzsEt8tSa/L
ev86IcHWA1gLd6evJrzCc/3+12dzCSc2DXTW28oSlTH4RqVa7qXydpSyPF2jkt/Sc9b5K+etNKLA
QMmBvOkaPzhd5kHvXmbNBRyusj0v7QkIOhS+MM7Tkp9zdjy0x50MwQsdOlsjiiuFQCGZ/VUOnUET
vKCIpalNyUvJUJsJ1MF8YlDdo28O4L8LV8zRixCbphtu22YkQDImtbscuIUt+m/TF1ygh8yfbysq
+6+GASWb25kPRqSBM8Znc9Or/0nn8IohqOW2uqMyN8QhsNAGeggsyaD5t85tA6jQSPR8BgAvJj2q
3uJU5spM1ctDPBWcK7RI2VCNgNsV5MQGrzkkmdPX65ihknLCsOIOZ+Cgnx5/3HUeBVWOrodZshpA
oh329XXr3lkeC2dHiG24Vw9SUqrStgfMGJp0fPZFry+Jgr5V+CuWgDaX1u3n2bAPa0bUvF7sMllN
/q3F4PnEMgyAoLN+qGC2Ogr0tlD/tgUE9sLk9nw/1OfDsXsrjiQtpG5EHq7y98scVm2PbFPAVh9y
wQJm0qzlxnRBN4zD12vd2LAZr3SlBSASZSFDmRywXt7Z+ZBQ51sE4h+UZFkz8VkaH1zAArvswqNS
lh4fI0avNGHM4uJaHVebqWPkohchJxKdFXUSjDW4DsJPgKUB+1CkxAZpl07vaUfCqDyLlwvYsmqn
AxHC4XYWhv+GncX3DU63Vi2V/S/fgVE9N8KmD0xlKyUv4iTZ7NSGH5/gbfGMMTaz0RIkCxo5yoRy
kTj6LyVzZM3UYDt2ku+Q0iRI6YwNXlEdjuk0WuGbAxYvfoF/8mr5fP95AdUbdNqGN34PmnUhljMk
tUy/azgdLDWJhIuMq3MpxKjcufWY1n4UX2ZQDuF73yBSJKGI4bf74f+dg+AY7R5Sie55dPoiD+xn
RC8ND7piPSuH94+ppmXBM+h0M6u0sViA1GUULTsDsZeCFrcZZu9RpPf42lF4yKuUpr5FUMs2U9BI
x2NRlqGtEsgCaqcNqIJy0wyZuDXaInxrf5z26iOh3Zb9+VW4X8Vyw/mg4NvbQxzLu/cHxAocF9BE
PAJXfR9Vf7ueBUI28CFgwz8tdapZy4g/KBIIYLHJT689iRqlT6abyaI2HCrGPJsyv/0l/qBo5JAU
Zxq67UhfJJhrsyNAIVRH1HUJRdY78i1O4ktdmjrNQrqrfqmsw4vZB5jyyEqWbtKnR6PsGkoj1dWw
jTafzspHKUNEqOTvH0+7KtTrVz2xITho/RyOjJtAKSSVX+FWjUC93aErn8Pj7FeNBB8D69sWymYH
5u2u266al8HuOegIpLkbMkF2UVmFl7ddCK2E3eM3XZV/iPrDN0PDxCnR/11qWCueCQCEcKvbaeRI
GfLBIdTcU6vSWKfrcrzGARYde2zU2XFpl/d4r0tXHLzEAwusGakO6y8XR1PAzsSezVi/LGLEnauQ
NDD+LrXYygs6zlDei6At/goAtzBWfjnlG6cFuMJ2J3PwEDL8uAWpTCXd/tEzPpUp+C01eLYfeOwJ
E3+nM+1ZQ7VJtB7VYs547G/6WRIDBaWxZ7zi6nMuaY3ob+BMSfKVToV44MgQmV+Zshy3bnfa3YdY
oSOu70mqToVKnjnanZ44xsCGIP+MESdc5lvqyH5SMw1zsQ5NPKkLrWl2FScuJ2LAx63uC5TTRo6c
k0nO4lqgVIWm14qG42sMg1B+C+g0v+wGFhtuDx/4R5bwuZM5JT5Kt9vrZ2/bwV7MZmXQ8BokV7JE
+djKZTdKUi0jk2Xq/vGrE9d4xRgc3tFdQIPfcYpNEKaqk6vmKJYn2VhGZbIhGYJ8F2Ag4G7UVofs
Ijp0pOwDvRMidGQ3bCGMun00NjOZT+aMvhufcoh4+9a9yQBIWvbKnncCs1fqVrdvBMT3U/R5eD8I
enbqi+taFPl7jdhQ5lNgiAE+D6LHiXxkPRyvQ1SmJiDWXyDbf9LDgr6/+GIG1HveSZsJJjpDU1Zs
EnO9kystfnWTuax1tefoeeIVl9J3JIpq8mTdm3OGlG+CQPGxRHlkPelmgwCSl9/V4JfckSL5QvO6
l+M6EprZvcz489A2wPRrLXfPAvfKSs3et8Fz3jbSG2DqGCNm3S/hALlR1oXvqNmauCyNUWfmybyC
yj1VBswjG9A8MODJWpG15SbXB9F+o1Osx8PvI5nMKiSMvdmGXmudHxPvcVKP7nN9V8oYd07PkIZL
8ckFtTl1m9sirpmXQj0UeTjEQa4hgdQdfzFujcs+z28P9wvOVdSzr+VbDqer95dmSvYhs7JQD3rt
weKIkc+/5iDsmfl0RsQIpedH9dzBk9pieNlDAYiEFCDeMpUJUQR4kHAa/rQ1A6pNQovGiLfFRYvc
tQpxHj3XqUZiph5gvman8sK3LiQgQ45s3AmVSvGH7ilI0wvZOpXqTAgq2xcF7I7hTWyBTJiIU+Fd
B7OSrLZmowNVHFw7sJSFKS6vgrvEsOrId6BmzR9QogBHVECwWILQ9WOmNQKK0RJj0SlVu15jdVC9
+sevqwtJBggKAR31hNfSNpgL7AR1cDDZRGL/zJyUd4ahEE8e2neaVV7008VDjnf5lHTMyqqSN9bS
FTZ1Ib38zakgLn1sgOzqSFVraeRvqrJ2XWlB/+JICIxoavBdbIanlOoMA5PxXWQLP31+VlP0utmp
LL1dRYQgdbWqpGUC2zBDjZAUCKQZdQcdQnOXjU76grPparc+7u+kuCOH6XFkL/hftkr84tjqSrL+
f+wh7rjXzBCKGbDpIPo4i3nE5iHc3pxZT3IVmjLyzlNQ5QOCaENm0/M2d0KsLoAw7S34acBm/vrx
Bt7OXbM7YcR9GhwYdQdMHWDUDqNBoY7NfeJX3NrP5mq1m0JxmemOJuJTNCjTqACMcDoJAX7TrvN9
xJ0CB2tVcWcx82bQjeOr8QfzpROjbucDlvB6AFDyeJ6/13nCvDyAH95Df4mMQwBSV+4lwFIftIRg
mzQsrgDy5PmAp5C7CbSe1CbVjjT98AoZsiSs3LmTeSD49F6ZqDJdqXzpLzv226tpNOIYs89gE0mc
CUdfLrX0r0DlH8HFrG5eVjm6HzCwT/R68WoU+9OQEmY92C4rK9skPenvzKZ2LFqtENbzheMKaz+d
YQjAgGbr8CGWGsaeVRk8/C5S8w9tct4MRPj0ojPFeK2y5Oj96A9xXdCy9g0cwV/HaIYJsO1/h8J6
r7NetLMfbQKt7RO3c3VnA0X2If1/CE5ASH+n3nuI06Yu0MbV3dfPWCAg2jzrWJPXm0VxpKI0vl9a
h2dfgsy2WCoIebaS9RF7FTkasbKlblePeWHIulM2voyGOh42MfuVHRZ2X9fJoa1FK9kWOmBBPVm6
wNzVD4AuMEM/Zwd3xEC1aMW49nD4sJ3vmgWWKOYcXqizyFbrbx7gBsqKPD7MFSeMrYpPfpw0hxwg
akxM9IeQ937FxqfToUJ67OpdxFjxh09K+gkv6t4HUErLNYbxXafpZ8O556umRAwFnb1ROSeOFMm5
x6vvg+rJ/WQJp9oe5YUDaLnyDq0P2FhCuOwHkUUTJotz6oOEW7PPegrq4BKquMk2T1e7TRWK9nSB
/qEfyFtOm1Tun1s50614kY4W5P2QPAgk8m7OBv844xgP6FiUSP7iEG+0VWhBl/TYBb/yR5Pnkk3q
62stFfxGUQJ0uc8GvEldfWR26oGmyv0PXNIE+DkIKCOsMYR9zG5ImYb0CEPvjuM909j8YWP44U3q
VMzVcmj/Tr3p/+vsVWANFYD5ZUeEE1vRUEbv3N43MKrZSgpNlRgb3i044rn2aMGChKZD7OlmAwta
H7FeAVNMGoiCn2aVnOfq9qQKxJ7+SmBST0JcdAsU3sADFCdlJRIzzkMubN5jMdBdsOp1OGoKe5g5
GA9w6g0NrhH9qf6LSi9BS0G1ObQQr/3hPZQmd8OZQadQPrsm/RBf0QXXkq3cTUZcDusOvd3ZXPqI
ZaO8JAbLLUoqY153I5meLSxn6bWpbeZSPMfBEmPuS/YSgtJmGHgTVFZ3lvF1gisTrgNmebe+uRIk
ZpyTv61bFIPVtx/GT82BOHvDbAZkYopdgebnHF8JNwrHYryjf1X9e5rwcCV5ccOIB+OANyfT377Q
sAzdlqQYirwuleK4ytUc2sYQIDHAi5E1MTCCnJufNu60J+owFMWH9vER3hrEVjsqjvzxufOk4fRX
m1JOiGdD5dQcNidhAdLjIOGPFer2BK5UzOELqURF1vRc9JUfZvpVcT/jmPSCJqYYpCAquCfLMwZh
ZFZqRJqPiDld18A0gxFFhoMZvz29aeD9hX0OsD+Ug1vidOcNdwSH3Q8IY8evKjojbu8Gv05EnP3G
0xFOOD1Z52F24dJSUlb30RPbtxsdFdjp+vtxTHQWNU4Y8FAGSZl+K5NxSTdER/IWZIHqci2OlrdV
nEjGm1boiMu/XwS7zYBJwrav/YSGzEIuTI7nXJnLTMBet+Rk8yJOh4tuSSQgAFXXAPUjPm23BE4p
bWLTVET2XqirJZ4B69kHoJFu5DRP1NaLmwdDP41iZb4KHMuDEE1oNs3LHIGFRTmAZJEcasiijyVI
kvG2RU2L6ksbrhoxaS4JzoKLR94r+wfnqTtHzAxWhWEPHebSq/j7J6m6Fj6Qs204zKVz7VQ4hcyz
qLtX2ZXVCeQQZB3lxQVdoogSP+X1TVNxqKqbBgg/Bf1AoMg9ZUW4PPRWjnUDK0Ck+ny9MHJvGmTD
+BoDxV97gJaoFoPYYj6vH8nfCKbCSr20nWD22ZR8b6rjfisQ4kMfPIYIco1Ef1fbcU7SjbHBEfDA
rk5WgrmXkcjBv6YOfXmLxvZxTCFNWwqh5rn0BV4mPABSlM4fDx/dCB6PFQoDcmDX/AzUxGxbY/2k
IfETAVTT5MSVxgOof9RMpi18cO0ikjtLZ3j09KLsisAx//IehLySVccgY9gfLBeX3w/y+bbGI7r+
4xKMxQXzEblmNS2chN8Q9+vrkV0UHU6xvV2VK17jBaL2hwvFNdjRy/C7H6XPT9m1rIDm0ybRtMWp
z8VESuIJlaUvGEXQ/skc/B19enGocbftKYpvqgk17UHKINHTlgfRMatCTVU2cu3uotDWubvAGvZG
l+aOLxTZB24QDj2x7AiA29t2kfEdF2WXtvOsySW8X5BydK3dV29ugSApulCKZSDwtHAZryZN1U4H
GnuJFFeZ7w62zNszIcCpxTomXU/Vz/6p527bH7ycSaHB70wcdyF6E1XEJGg1iH/P/LJTZ4bR8Y05
2GU10Ay/XNTsRJYqyKXqj6rBJHH1v3jPHOwofBdD7hOWwfaSAbnwoFGlAy85BJgH7bFnUh1DcBuA
9nj+/YpTSPFZoQWQEFwLLXHnYdELPa8Ra/M2V6ifDLwvgYhtIdrRWh5I6fGDNdkD3zu7UVdB6t2u
kTFySwVc2S5CrB2geOQ5ZCpuBNbmuNDteC9S1A3gLnwHr32BYVGj+KJ1Tbt4oXIfvp8KHypVyeBb
N+7+vCVFYEPs5EffMUYOBJ2+aacDUooaznK/KRT54e0Tews6E+QKUAyVdrIJntBN65SiK2CZjDCI
YVcoeUzU2v5dQDiYSWXCp/iryNmwbTWz+92R5dFZk69dMRi98FJJs4dJWZDm6uEdIq3TgMAkE8/4
pjy/RQFf2hx/lNgLOmaUQ9O0YnziD4hhglappaYtT1I6nmssZQMrfOq8c/1g3FB32dZCf4GBHpuB
2ene5B88NQXbOJZ+V+HXhmNb3DEg3emBuhPxQdQG93aBLxV5GdUtPiDT/zkyAa8QYLxOqbBeY7JC
ybVaculupULM+HxLpTnfB8sGIrPkzF3Z7BZX1XweJUGvbJ8fWCSoXFI+6PG4m3TkQt584sJEDpNI
pNFTNuPuzy7/mWthCwonMyYg7TA09YTyVOy3Lkw/3UAvf74G+CzUVgY/mnidkmD7uNtYpHNCO1Pn
BEUjehFGPpP2i2G9WQWvvo2jnAHjVeLcY4A809SkihKa54HwwtpkC4OSmZKn0tG4AV8soZ44xBoM
R3DzjdRmRq4AtU/xL1TVh8M8UPcMVn+9jbyhwqzmAeSbvFBLl44KEMQnNeIg6Hp+mREftfJBEmp8
aiJDnfEd2pb4dYZSWgfTCmJoI+ZSRHDxCCDEc4BQ49ZucpljbPJJsAIyTRz7fgXC4o5b9QStWjWs
XF1Va6H3+I2QaUEYDIkezXpnlFlCA/NaAwQ3sfA7TXxz9JPmcVgIzO8kNX664LuPHddlcm4KnyMI
hhhd6Y0aywzM2QYyyvPWKX40zQcMfapHVNPyjyk8/iATeWNAFeIjwceC4eiG1N7AWq2uquFuZkyR
H57G+SnxhIZY6fAp1g7vvUiVInYuckKwrwUCTsNiHriclB1bUjSbtlYVWs0hfUZTQEw9ne9C5mBp
Fp9AdMn5o3LVqezlqXZnXN4y9k0hrrayNiyn1lJooLrB4albMRI1yEm5t+bP1rTrHfETYfnre0U5
tNpWH3caHxFhVQ6L1egRnpuaMZ8NlehFQHT9lMcjIfsv9yd2X6b3DOV4y52x+yUl2NaeRZmmfIeZ
Xtlh+sEc23qvZYXTO6dM9Cobk1rQmFp/7i9uNc5fiS2MLBv3dvE3Yv6tt/AlKKl+5gbeymyyJGR8
yOtVnqc5g5/P4lh3xr6nf7iMxIefJdcEv9RU1XjOj9NBcq9PEEgo3V1wAW5kXqDAvYS7AzUxqp8f
PuzVj1cNCad0qlcotMz1f6HclzZMXKTQOd4hK4ilBvpsHSa15HmMYpxa446/ARQTBU2vigpp5znY
uQb6zYlNRwZ6MaXyHfov5mgCKDsT+DPN7EfYkkklM//hFy6PewLWggHNQmaCzx31sziaI7rM3PAX
TbBoH9EsBEPYK5KtxuTC7tamITkRub2wdlqFjMuwz2mU90hT7r8zDjj1VNulrIy3h6EWmLkaAEVn
6efpPs2/oeKHOvdZN6BikMz3hlxWONkbIdMWOvCf5XQGAm6bCG93emF5+SZllB6AQkw/G8qGtXW1
kFKct7bfEC4OniexaFsg4v24njSai0q1wQUjcu31Bil1774UGHZ0DRjOSKihH89zNmm+vlQxtGVw
ipffwUZ8WcHbaJat9l4f8QTI+/eoiro2owQ9GjKcMOQiKeJzUPGemUd6bxNoGfWoBjt+L0AaVqkg
db0tylFu2CJok/HM50fyg3ArMYht72a2pX/xszlM6JMozv6XzI94E91DxRQ3LHLHmXFrFjvDCAMV
jC0xAoUCy9JpBeUVhdcbXzEgeY6U1trZyL0vXdBrP+jGoP6Xo+N70Na5ct3rlds3syzPwIClIdkP
3z6IUuqPBBc6l+7CahfwfzdMMcN2prpZqspMAD/a34D0IAy02taksgTvGRbGW2m0RKLh0N7jjVry
F6oCg+7cV1xRRJ4j7eDff6shlbr2cieurqItm8zAqxzQjpdfd6G3Pt7+3ASiMkLh4cx6IGNOnuts
LSeuVpEpN900QQXDZE2P7Js7VfDvD0GRvTsjB0wHz2vaBsJcdsF65vlOHf75OFLmrMPgH+KMh2zW
0c2NN6ka0BxTSEl9F7rNRtYvAw0bc+b+9WgL6MDY/FN00UYI8O/kquVPfjNMLv1FiVHHvUUPu3n0
6IzbTDAtXLMbIomLoj7ihYCbEXAd4cAd2OVBchYuH08uBzEyc697wWqgN8vrhZ+L+KSiaK11tifI
iJXhLMfchfnijznjStapTEtte6dIlvUfZXYQhlaRhJuxDHj5msR4CVaSD6FHKYZLjc7M9o9ZBkbe
/KUF5Znqkf0i/GHz/HILptfhq8Vm790jT2zpOlFtSPNHknVX1eWLlXrDaPqne9MD121rkmdRFb5S
lfqsEQ4wTmAaDbarAsIPZSSogtyFWsd38mAibXca/Ej206AzNLaptoBqae/HDIK4encWFBuaXVb7
wGricVCpTpGwucO0YSbH2Bu44mspIdRDpH2yvriVx1FmEgq5uN4y2xMqDcs9r8fv4iYS+ILopU1m
WDk1ugNVnP20auM/49LK6MLZRmm9OyMIm8uCMJvjzedhLB1Pg5k4jEpbHPYuXQbQ1vLwE2Z2M5OS
DDm2buPKgXoZWE/86iywrtaDTGpnsLQG2DtHTLoi7xfyrjL1PboGsykhjNp6HxsCSE565StYXaK2
pZb3U0eQAvXpVUfvyelbw0gaUPWDz/Ocb66eFFtz4MgUN0jeJYnKk5XB1hbQvcmW7FD1C8cA8zay
U6sq76xZOAV6Iakw+8An9yaJilhPuncGCVkGW37Y6OH8z2GHnYBMO5+xMRHgMw0pmZcsdw72Vj6h
9qXQ9CwmwBvhTKyf70TDry5fXQzoQeKRVV4Rcs9xrUmreCafMosE5DG/qCbakxpFVAhOlzQYzJhO
dd2jw+J5N+h9CfYMczCxBExachaR3ZsQ6aBxCYMELOqcoCEx4xVFencMzkeL1Sy/SNSKKhSimagu
WtYyNXNIYTGvdjBBW7OJtR2dF7qtm1VAxLQA+gaEPDF1BV86GATc/BYXUD/Ihuibd8Wy506F95Jy
zs4MRd4sUyXj1ik3ZQusZT8+8A4vG1Txs4PlGuKdtnF9T+uvAXolqG3Gfxge5lJUnrJSUvNZzpGa
g24tqJwozITDU2Dk3fhaUphWQB1YhRi82ervz1RgrG/hFIKRgpkxRwwlcLETpOK1Ba71dLzNFcmF
TG5Vu8/X7Qb8FzS6xgSarjAyLtiCWukvaBMN+sG0lTyA/Rgu002x7pg/GOy1RsY4dGB92V6W037K
i5HfTMlVOlnGJfYS55knacuRmI0OwJgM2ULqHN9LymqFvUg6dTa4xQ9Vg3pSz7mzpin290PMrhdd
bCZFeq8Eg5wYQ/rACcOCtBa5ez9VI1q1QvBz12jeAZ0b4bSKHZ943yS8729wffeXDIDTtDxk6rOw
1ZT8Fs4l4FsPT+IBqbynAOJxv8foYGErHsnaPMwwbvqeHmOKirR49v6J7B+6MnZth8+zP4Eb03xv
Y6ZPE/vxVFEmFi8oOEWKe6IJ9sjth5tynmih78CZxs2EtKqMfSnORxMfQe/sQje/aq0PV5jufpKj
nb1OAeVWAlS81pvA4P8twTTIigab2VIE724WY11BeN2k2omv87zRtwuEfK7FleVtNvslNPzuSG61
jimh0MkJkFUsOljg0YyRahvS8h10iJHweIL7aWN0hmigtLw09cXCr/ZyK3jUMZf6kNXeew4QDkVI
e6BjrbDtMAdXGwUzw/b9M8qS0io5YXPgQDhaCW9BSgxXaEkRbMSa3lWlm1XpSAHp+LjDQ/4dChXH
u8L9aHV3y+Nu7Z3BTNKQ7r2DFddhRsXEfnFNeOvSw1q8L41xVdAyCJni06+l4TrvjsgnJXT/F/YM
8KTOykffbRoi4sD+VVHAov6oybXyQNsWaFvUf5ZyIr5jOwr5kwMaNZv2qmZaX1d2nZfJBuSd/KCY
KTSxyOUJnmwxUMVDYA4o/8NWEbyEABrKho7XdJHhmDrvVt2bt9WTR0rIyh2Bn46EuJ3owyhD+pva
rRgnAemtLqUW7mZevDnwrSnVYgq/MnYK0rN0N3laHIEg9H4yMXrWB1LNQ6qoaOM9mPwnkUSO3ys/
MHiulkqNY/wGQq5uUjyd3vtocwyI3Iezbvr6HcJPNNwS5sUALF/eABrn/ohXUIwcfKl3uTXmdcb4
x1Lph6aKycFft870sdvsv8dGDPNo16pKQWoHbgCsV93JhRlILja1Sjis8NbtSluErDn3Br+MuVLm
5k6OlZcZfsQrsQM0jh9pK8P8Mge85obE6i00GJ3S/CHJUlH1xfu7WR8RjB/bfS7ye02WQkvgW0X5
HgnoRmaXpFmjv8ikZx3vp7B9bitaaPlTkySZVOO5TFwRRvYNHSfwd3htax6DEiJIUS5YNluSM6S/
faV0q71l6B5BDLNv5jIMaODlEvWTflJzZpXLKZQsyiYPrqJlp0Q/0527H+IkUxfFQvaQ1/UAnPyJ
FBwAYdgrq/0d1J0XUpvxryTvwCe0FGldt6rN5CRt/OtN3w2ULmAXStEMfas8ypdJdU5DR4FywXug
fPdrsT5YktBp4sqtNxRx1B8yJrYuw4Y8JV/7ztiSkJffE7XZQbW5fjv+RbDtRuXWTMf0KilNQfSr
oJgkK1OlEG0mGZBgb0XUdTlzYWfO7chYWA0/ekaW9/fwISEfzEhYSlm+5LvSk68KtABw/SWnLAtN
554iEpLwQIUBGsYQ5TVo2/66/5G8w+RMiwm4nqWa3p/nBMa3WCjzsjxySrH1BmaMgl/qChhl+dm/
MYp5LqZJKS2B5Si9h9oYxGU/0QU27TpBwJQX9yx0oF7RFE5F8i/sIU2mMBxOeAKW4MgyizJ+KFaZ
OVGXsSNa7pkcicBK0u+NnJa0nQ8z+0O9PpmA4oUXWg35axC+QwuTs12kf4XHqFdFpqtFZvPKjsvZ
U0Y8lkuZ9xA/hpWijllLevOxKLg5p0H2QPxFcCGFXETib0/s/EqDTp3GNQxY8m0E8xAEM8ly8kYg
ZqUW9IsOGG9n8j3uHjkf+tADN4i6S47TEW7q7zAHc5fGIHTKiriu6RBe/Bw3gGqYFk4nu+vz2ALX
irJTVbqVgmid3Fx71h2F/IU6VjLZSijOCFh5fjdId7tNa5EQFRxR54g5L+tgoLriqRJZznN12/qb
sTh4fl0UDqTWHpNcD6amBBB1f0wPgaJC3dYWxjO8T39yvQI/WCXjz2nYj52FRIKMQLn7hHY+QFef
NZRyhdZ7LI8xplJJwK+7oyZAQfUkAsrWtEGQc9j+lMgqaWqVAiIZf6KnINeHHoZDeJaAa4wv8zKr
3PHTq2yyrexy2CDt8xHegOO+p+ltBqWqLrzt1SyIFTM2j7g7DWMdQoDMAQJpALsUXEpVWDIOmIow
0U2GNzn6Awr8R9jJbedgdKappoblM+hp5t5tTKrV3uFbIVfufUTYxPbAoyye0M/59zDlCGqu1QhL
+CcFL1AcZcnpdrz7I+GzULidvzeovZRre9ZyKhf0WgO+Ho1J3rNbPyxvs/FH90vMjmTF7YYQRfIE
Gi4ZD6Pm7Ej61Wutkg/M3yrxlty/XV7nNjFC880O39n20oaUjg76VmPjmJYC828qEFy2he9dvq75
Ncv+piBgYHh+vx6TGUZkixvFQmwuaLIDczydZr0LwF4dmwFUS0819t96x0zzzEdIG0uwrNZSm92t
blvkb2YugLz6O+zzBkvIknKMfovjy+PKMpGZYlMTZknCB7oM5EvgHg2NpP/owhjgwyPXkIS7NHu4
+/+Y2+D8UnWc7kuUUCdcZiqBQIsE/kH7NRYMu3eaFbB5UdhWfSf6syCTD2QxNurDs58KuLiobUs/
F2Q2LGPp981c/TQH52lOQQ5ibNAlL4ERHPbdhnb+21Y8Ybd1v9Xml/YHIBCcpgriKL+4kwOSzgUq
miW0rgmqDz70K4hcKwB4oYtrRBsZjz5mSSUgKjWqt4RRzlVK6r7PH6wy/kwIa3BxnOFukkZuc5c3
K4YBsJWYzzD8fWhh+t9K3aBRabS4mLvaToWhOekI9Dg3MDEde93BDOlEJN4sk2UA34HFffv839MZ
LwkimxxViphD2uZ9qnJ1kwUDT2O7sf9gPtasDjNaRqfHsdn1dAyqXJ8JYE2cx7LSNieEbY20wn85
FDDmpUnoueMb7jI4RACzbTcUfyINpYzHMVTvpNSgsSimKSPickzs83d9hVOuvZB/XOqMNdJwsfZ6
kaRj+4AnEXelpIM8KasdyGAyohdtMghhFzW2q08AsgQZODrQP08GqHTCyOHJtj2c0F1gbQuNyqaY
Bp2it9mXPylfAI/0BeEHcmFkJvi5R3jABA1GVfZ3kLgoGExkq8/EKR9cA2L8HyBR8qFYFAPbRWyc
4xoOWFNrp2U6MzXyPIXa+qp+8c/Ts8ZngbynAJxjzmfQDhkDyl0Pa2bAPGUvkduOIbGhkhA/OhW7
d/METTuNdN2i+hoQcB1egdjNSw0mRzv5hjWsyOKdVOgz8NC1BfRBC5o8/D8QmfWFvcZVmcVFWZ9q
+WY70mgI+S6tIbLuQyFoMD2bgK7g7k1aGvKfzzQPBMPG367o8cFn4BAvMiPqObYlYCwvdPRgjyEY
lIX0g5NIc/9Tivwb85TUoE51rRiXG3EBYiLhytxIQUboE+pLNwEq/C2HyoB+51EU9uuadpSP3M2W
EApbJKWmf7e5Me9Y94q2qiXmnhuB5YOiB5feUYmTD03z9eO0a/Z24NLUIKK05xV17kqQXEyqiIFA
4VqlnH+TuVPQgC7G0LpfYtssIkb8u25MzDc5hClRbFUdT69NpJOLp5ynapAxYF2I0feUr6L3lWAh
vcdGQqwI5hvrY89cL0wxyNIaMqhP97dlRxxFc90z708YEKXYc59tQnQA+Tlt0QWxTCXr5DWHbF24
EIL2qSkT0ZwtGbsMyyzaMGwC1E1LmK9+MlnowAhkTOJE/JTtOdgDD+xOAoesL3kD+b7f2sonJvcs
m/xPxnPAzGPpn+mibPr5Gsf0AKFtcYcoyX8jj6ytshAIjE/KB/cGVMmYV48BtGC1hMwDM5PYqs2f
yvtHzK1Y7nsHTUU9AlohlCGxnNQmOuwlmo2atjo1shn+ogHEi2NU1nZJ1sUWYII+8IdfPjlHM47D
19ettXN+oXvwwu1ydfIxXig8ytfzNbc3wtY8p2EgKTQbQKmgnEUZ/ob2U47sVPafgD5vyK2hINgA
7dbQ7OdLlJONqyz5H6EYYOz8Xkn8N8yFLtY6/9qa9ujZW99UK72ieHnsrFdljy7SCfXewGVr/y7b
tDHB7Y1qmtSG3aguR4msO/OJXfBzYIcTU+dKvYViJmh6GESNWGimfKYqxohWmWVMnhhm3S4YTL75
BobgegjUxoibTQXB1EDA2R4AJQsfqgBL1IuUFdkMFyYH14XMXfgzT4AdVUKtx3Y2jN6o8tBaDeSQ
DOkBxmggZSG0NTbRXxbev67pA969Kl4FHMBtSovlJKFyNTghqM7o0LQGOvWqcF1qr6FZ3CgQtLEX
W9sSnXo0/lB3sdjDLBzBijRgnbLlBpmLHFcICw1lgXMy02MwSpdKrS6ZJdWduih9eqE+sP2vnYn4
vUj33tDW8NlhPMVVH3xgyfmfuqyHlkAxlThQA1woF1ensxMzMnNCsSl7nf1kuPHcQU9Fy5Ixjo3h
NPGMrTd+nHcaS1fMMUJB0xFHPXJbRWqiUVmqqBlsQ+XhHlbruRPoUQ0fX5QeM1DAaJs3jElxYR+V
meNrHvcvROQQdRM19cdH73Mye60nLMcgOi5Ty6sVawxVRpbXC2rYdKkFMpZMPECijLIdGoIfFd4d
JhuLpP9GUbXuFXv67abjbS+BqVU9K8voAM4f1QOwb9AkPi1ogGa/ngzK7fTQFaEbTr/KDJSAO5Km
E6iX6xlOMmXBy2qsUjzhlYU9z6pou9Dl82Z/GEKzyMXgCC/sBrlffEgHSL768XQHKyTBg3eVuc60
vbsU47UM/WtLauM6oj3hfMAm2uHCMccmIN4YY8QNYHcQsht7JOcLOBSPYmGS4yS4rLPTX4rDA+aI
l3ZCkKJr/NbTJNNOnFgMZBpsx71fUw54IXVsecK5r1YynANFgeCUrivZb0onbce0Qac7HbfM1qwL
J0CQ9wqY5GA+/y7SOp7JwFvyH8f0FMt4gZFDTLuTn6lbV2jIBKgDtyQrGV33JezBf6p9jTi8mNti
nVdC5869/h7PvQL+Z3TEE4+oaTJBprYHvZ6RIZE/Tgj+Zeh7hW8S8LLB/0NoxhMBC47jw1tc5bbC
zx4xT/AHS5XzfyEFmIVkBFpSn2P8jHgJpA0vfBliObSsxdLhA6TzrPyGn7km7bT3fo1goJxzj8YL
MSOQrTaqvyuk2q3Or9D3CGmAUiO3UVL+NYnkeMxlahB3FhsNHnzS7E3hpVJCMIudIvZtvUluzNzK
+QXGho71cu0rZbkDU+b5yOCnpts+XmqFX12TzaBIuPh6kHKems6c4saVf8O+9xoWwyF9Ga20KDjv
WOFeCuDr2ZaJi+QpkdWzKRoqH6O2rZd/KAncmeaQRWI2E8re1FcvupCwIe7N9xsONzlXFicqnPvt
U7xt4Kg9xWK2tJxM/7FSr1BtBo2U3cY5bFl7QNT0hzLGVMwl0V4aLreqNIbHp8HXXOULwY+JozUw
bn0mngLUPrqOsn+ltK1n+AG5JOoSzzimFXo/sl+8MruXeNu+j/PqfIDi4OJMrxtvmfJed64bnDmJ
bH6RNvJrnHYzeJxnFlaR8hnUc891asFTdoOY/9rX+kopGOHKKQEt6gNRfhYEWVf4TcbBfRNJb9xO
deky+rL/tN5UJXIKVADhzrYCh/MI4ItNxKO4bmDUnaGSuwA/k1JAjXHnKxhPStqDDrgUAtsv3K0Y
U+fJ2oQr6j8/061jDBSppMiOmEsQdmGsx1fkLIBlfoWERn01nPU0pgSqv5hCU+DTFxte/DUEqMma
8axyhhG4jetAEj6TkQZ3ptNng6KJMaSxEodxyH8x8aG5U+wqRk/XL2ZpLdP/r7Yzb/x/jLC/H+6N
ZwqMYOprhRMuhUSzW7f4/KnXDjOs1yOOAJ2aWpKoWLybzZOhtTWpCY1LN+hkPk6XB16hYovuywHg
B6YCOHN4+1irH84pkddGKXwPgme1X9tIbZFhvJBve8AvWZoudER5rEGChJ8Rwd7v9dNf0Cb5Dxtq
uOe3ecFwLNkV7e3GyP3xyqMUiLTuo/s6WKBMB/pzz0V8wMdyYG5W0XaQHijwkGa2rUV/QzaucPOV
+ZlENGCcD1Ty61VqknfTnfJUF1G79JsbWXA39ylnjGwKtbdky9QILv7G3E5WXvtdKU22TIqZwLmL
zaaOirGwNWmimU/9To4Q7TernTNarhzxOKP6cGemjwvqUAwsSgraJUB0cBIqOA97mbHF12AEyjeh
AiZ5wcPewFkjNIFkzNIf33uNpRhTNhb46DuhpwLZ81dFcPdhmkFNt02qdUQCSy/KATGVuSrVXPFE
UcuHt4rimimW9MRpHoWK0vDxCe3bbeSC4eKFS14xoFEPRNFyK9KW88zx1jMZsd/it0vfE/bP4AA6
k4laLHo9mCkv+/LLPdQFkFy3g/dRi1DqoM701o3YUJitOgY2UO1bV0dyYGVku/wSia3pUfwgcmW+
BwPfLakaRFf0wFE/y4/+ZuY9nsMdo4NrCF6gLTge7M9wSp+mos/qr+mA3zCnJIcgBxRb15qkbhQX
LCP7jODApdE7Ow+hxJACP8i3z6j7I34NE6MFK8WwpcbxgXHWbtwYiLbjZtByEQHC3Ke4Q//FaCru
aq02n9Tfvkfd9vYPfoIzKm4SMi+vi+y/8ObpLBfIcrEiW/QpQDUSHx+CRrK/SAV7B9i+oLghUemC
uktwUug8e/2q2SzOl3mJONxovdn1zt4sJ9vL/W0eOdTjKwPiFgMAcB1vd9sVmv8QBWprWojffS8P
nqtJUq3VUdNjmUuKv6BLzfMmyUY/WGUTVxjMI3ZGoriepvskxrb/bwqGcGID4yTWSQaeymr2lZ97
YR7KH22/7k131CpoDPdOMvx3ZioMAxEDO2pt5vruHgsYRDoqa2AkHubL4BSqLSb7gdyYcoY+iC9V
DAw0R4Gd4zI8l399qNiWpXwhmwfpVruVNdIDE0SFjZ5IxT91KLNZxsXDYx4GNrYcRpUX6AhvQa73
lMnlTeOv0aBg1A3RDIVNRSgrwAXmPWSOvto5PPuuFWeOlwEAj1nb7kOUDky1quEgnWD/T0cJu8Qt
/Ehpy2+t2rUnmaN4gbQLL8GdjSLdz4b7EdTtq7k7SuhTkCLsm4R9GcaNZ2liXXKfTak/e9WrbWQr
xXtR+MFCyk2/jCXUuJWFEyAcyG7GwcSzLV+m/2Aeg3bfiEIS571INw6d2Tf15dC0aE8PDgpJTEcT
9pUCPYc1SVEkRz22UryFiKGn+ecstQXBMLZUCwL8RSAHBu+InGZ4SeiDI6S1v2eIIPyIxTnGWncc
iGdiJZFDA0CkcjKf5GJeONNIKLtbM7Gx+E0nfndH2K5sVjwyoWMaYkYIgWuCKySFok9VXYG0ngCf
Xsfz+Occ2PTS+KlJXEKj0Pu5BEcZoj0SuBbVQFcqQxi7DCLrkGqe9YTj+4O/F4r7mo9UxxsMNVya
hHo3lCgsre4RVA/8DS71/YQ38t2eNZJ+Igh1Xn5+/8h/Uxtw+B6m4QXuZjFGV3ijHJZZBAwraL98
ARtdwNSsOVldZEtQL+hxwj2DDuugd8DLw8WS8R7g4F5UBZ4I1LTiTuZAy1hytBcRYhR7QhnbEYdR
BkAWH6ssParoXcGsSaXesOjWMn+ESNIp79aXyi1tfuFG7R67etw+kvDosf1ugTx+Qibhz5I3tpWY
oCFFK3Y9XTxrWNb71w9OofocLK9xXQURtYGuZRtuvcf9w+R2zrQhM8meM4IIsQUzDb4b6UXZSxyZ
vgXzHuUukDEAAi0tSHvb0H0LLiO5Ya8qQ/aS6XrvkavvAtqxi1AmCr5SiXF7YFOU+k3SGuYeyM6P
94dNhmmkNROgn9W3/Wi6Cf73e+/CcRXS7otl8L1ha16f5XyhyE6n4x5/bZ7WRC/E/DCcBt7JtGK5
AxPWqzuWqomKtxD8PpHWWgs9pSxvb0WLxCO8+Ps9eigw/AZgouoh9U2KGoy/F/2i7Wbzq+9rCCFz
9E+IcnKnUHVsrjlwY9jVSt1xd4aJcBTKSa4oqzRyJ0xJb2W/XYRHzfD5sN7pL24TStsao1dbhXlY
iiL//xuM0wYmxHlitJwymh3JT9PhlGvli9DOkov8ewjyPLmm0iPlfSitZq1L6cGkxwsqwzsIKW/Q
gP7uQTJIgIimMQBavUeJyR3POzkWGMHgAbiZvGBeTL1LGHuQjpy1ly/5AfVS37tlat8tsykH2x/K
42/1LklYYDzKPymcPQY66Eu26O2BEw6+ItuWlzMxI8Q7J9rGQEnl68oaMNKKY1qrv53UiRtiHcWt
5i2UmQY3+Fp3TpbuIAuiRsSbWiCxCd6NCxFvAV3JsuHpV4g0G5etwrQ7lW9KVooMYzWPQyj/E6UW
y+/rwBMd0fWqmq/3ts4mwq6QWZYuyp5TszM4p5A5I36losBoSU6SPfySNaArHWEyI8X3CQTMlJWq
tbYLMPzoLpRL/rWU2Pk5sC2MWaHadoihE8vAE4HqIo3sXy7O+C9D9ZziF0nZGa+kXiQgFv0soiVB
MTr0Ietn6U7gmqAWbYR6nt9U5MUr/IyVm7V8aNBAfUGzNo7Gk0k6tS4dJaURBrnPD9Z0+JKgPspL
AkMww060BapkIVY2VWYFME4Jtf07ETF2jrKbyH/1uLTureTRdZG9FxuCEk2Op7MdnQQRvsKW8z3b
iRz9Nlxux7RHN500S46zYb9H45sEvJWt8DMBy0+UnF0NzTRcZjjMeTM9fOM4onHXT5lWRJeIe7XS
i4jRDosWWDlEh/bJvkQ13qJqAEpJjurOuVIB9z2fRHz8CuQAHW2C4xFr+FcYYOqqxK+zfQcExdCx
zCX5nbgknTVDhcfwmrlyRKCnrExo47JjJECz0MyY2NUE1DH8TWQIKiFLNfuV48kUc/EcukK5unS2
tbSc0Ptx4M4M831VH82vCi7oXZVqezlaAGAbigNOcICb9l8u+DZQD8BLFPOXOPZ986uH1D/Dw5Or
O07b/CCsLwhwaWdYNARTU15BUsYO6Wfij7lBSYH6LwAQExbR4rCK0xs2f/2UkONIPrY7iIFn/cSQ
KV6wErXMBANAE089flZH7aqyKLgv+yykLopaGES66YFc25aY3hgf4aSGgdq4qWizFw4W8DYOf3MO
HFxQRUmjjuOPcH0Psr+pR6IS6tMUy4ctXBK36Njo/LY72xiExibgbhpxLCuidk7T7S58PFQLrc9F
Dm3y79M+vnwuurnTr01S2INQFYdaTCuOByEN/SwITz6f+V4rv0iDGxgpKsKWLzP2/HvEGgZHaK+H
JzgfSRy/a0vaosJ7i4vQTPCUKlHSZhLP5uujOdZGkpm2C76/mCKPECzphMURh8jyVI1+wBnYAKA2
1gF/Q37Kk8X0AJgOZRwMeZKKoCLqoBTjKzODPatiieeNyxe+W8Fb3aKYFxZvPyryAP/p8ilUIOwy
N5GdF7dExR5lLnZNB/ReZwVgdcBPSlWcZi50psxfL7DfZciETVCafe1p9OQxIlGpK7aKTITSxRD5
WsX7kr4lbu5pXr+FyGOGq9bCD65lFv4d9WYjxbsLyu/J5A3jb/VasJ36E9fZh3aFWDCd02543AV2
1bXk688omKq7+n7aqcpQ7MRCrpwDK0gBPq7F1wWC1/3jP88uXwjJW+0E6aEVvVpVENs7BHmN04Ck
Vuasy0GmG2FXA0PQlv9oMF8JD6KopDv6+jcBYK9UiHvX0DR6eeKmcSKLsfs/AbzoS53ad5tJzCID
f6Ns5qRrNtw+pJZjL3QvaBH0cO/04goS+v9qkZk9U8f+wedoCD+K3zx3pqYXOWvmjHk4Bs5QVRuV
+SOw8lk7IY+G1kNJdiTqLnfValOlzDxxQHqUeqSB37tbLG0mMrN7pVAxjfoVjP4QGnGfh70G1GyB
Cxl33gIEQhH/3Yhw6f8aO0Szw89pF5Yca7YlCaa/tZuV4XRPCSnrPrch7Pue3ma9wXp+Hy/2vzf7
wgynQlxmH5zz00j0fuW/N7YNWu6HAFxVyVS9FyTNb5oy3YE8WRGhoZ24GoKkOt5Ecb1QjtxGY90R
9ClP+fTMQIGePfIIo1X0hfCeUxRP5SFKqHplNcNzVkMTbI89WLqBBPgftlHZPoIScuWbCGv8FykR
cST2aVFa0TceLbJVBnrBQeIHsq8ffbhvMa9XDo5aOQFlXSs2hJYudvINqyqHVqxG9CDgilmbuPJ+
05XyeAwyPY49lgV3RltUzy2+7DGE13Bk5Ulod7DoYRaFsOWV0Hrt29lL6CpLQQ5wSw0/cam/QwhO
Ni1j6z22BBgTfDfr9rBy/UJJO19QD+Bnw5Cm2UPd2ACGTlqWSDYMBzM2ZybLN6idxiVUIFG/eYqZ
TjayLi5pnX9+FjQ+ePzVHF93UjaVqcMkykERGLC1dfX2UWbSEm7lDJuVZL5t3EtY88/rgL8iISfz
Nv89nRfDjaAgIoM4D5/sQ0I3n1zR7VQYBIrHWBLVoOvWOEE+5AfuBYxi7mGLzFC8r84tknrQsOVV
9aQ3m0q2VNaM0Kgs1rqaLNKa3A+3MflkXbGdFUorXNarGOOdRLeY65xfH2afD5Vt99vsj8lpS2D3
GH8VZtLowp+11EPLXatD6RFh62gPVv5Dy/UsKLw1DAaXJKgbsCnBxEppFZW0ZNEcX8CDEMaRGcon
2R1Dq2pKdkNvN4bihGguN3wdjndti6NLu92Tvs30wBTBcpAZUyP3fOa4l1ccWByqtyR5ynouZGWx
i+F5oivH8J14d0Ajk6V7hPBGLobeRK8SuaaB23ij4tAV/JdoQnuIqKft/A+f3JjQSdJEfPZ3otxA
pId3aN4rQqI92ysSlvWIBJbOojJIT7gzOQlCY8+1/toi4TFXGMefRq1FKAaDc/OvevABQvdRxKFA
vRvUxE2V/iklNMDPKaACetSFj8wN9V2SNg+XjvJTsVLKL35fAH2NBqX1M4E96+odbAzuAxZ0KMg6
sKnZGFVanm1OREpBlCeL3HBG811IpnOCBrgJKPzaeiosIZCj8PIShiGVG1YePbuc1c6DsIAXoFzQ
bRPTKaNJzM9A3vX+tdWWRtNN7EJFZOPTUJH21YeKbjlU1VdwzhXN0pyTEDjl02a4wwa5x088aL0G
f/k8cewMQLqBK3J9RVDPC61HGNOmatVRLbdInXNEEH3WrwBmYQBo/XaSJsGu5+//zil0mUV3jSbM
J6v4olWbHY/AqzdPm/FSemd9onHFgCi112OJjDNtQs8jVNojq/epFhpsVXryYRyGG9uVIAxcIw9E
LRFZsCumOUkmJp7HljEuGnbigiNT+OwgVT/2oWuaY/6VUo14dlrIqHKbeHgwj6o6F8YIkka7qXm8
BoYLWoHMbJfuGdYQo73VIwaB5Gqa3HtejCg+vwIZgvH0tJnoU+A10Km4lHKQeu2k29VJc/Y9vLml
TutdGZq9lTaRtGDEvPVmMqL/9Th/uW2Du9jfhD/MG+nUlkvxp+dXwCG26YYGcQV0mSfaQ3+k6z2g
AVLGY9eSj1hiSv25VyXjBsahZaBG1eQg7qfnFr5dz4JSN415AbXiRDgu5HRdulW0U9Bthp6JXFx6
PeYVq8mIsMIN0dUc+ldvDdUPwvZRQzXYsy2QSf1cdwMapwzBdcbcWdHoG/9wbuhypKAhETqOz1TI
KZ4Y6BYJKt2lmmFcDnqsDjyRWvgI8CG0Jv69ctysrfBkk+fZCkSV34IIatkY1fNJwr87ekjyL//f
qqa1978yaK0t54Z4MuwvzNAgAg8/gh01+kqPeRX/mpLbQ0HIF+gSVsFEWdL7hn5FAiXlBN1mfqWo
8fvE29x6SiF1lO5AGKGufo9KUeVbj9TTWzwRjSB4Ee0rDjSMMbMRAXMx9lvc6VN6C71M5fjan4FF
LeTJxUKlu58hFmD2dh8Dpd+Dr/vSNgMIpFAV80NVTY1Ite8roZQVhhBzQvlREHkQafmcAAFbqVLp
oK0+v1WNI3r3Ql4uNkHiP/oYobyAXLcGjaC3VyOgbsPmWGHPu+rlHB6IUuwcTeOnoJaoFu/hgYBL
h+f9HllGNdZUQVGJye6ZZ3FXoCI3pvdk8i1Bal08pJNzhFkioSJ0+/PR+IJ+gCIBP4WHntcqagE/
21pCJsL92TLd3ikdgFrrwOxe+ZF16XuoaTrswtvwtm6aIuXc+9fRPwPbzDJ5xu//3lQP1aGIrGsK
tpH80f4xlwkyRYV4IxcZNGaGPeFrSVkz7lk4BVZBySc7l6If/TeQVfeO5J1gJ7HnFeLH+LCOmPs9
V52dRuab8H55xPkM6Zl1LOnvMYVea/d7fuQIaEAMzU1ZMWMTZsZDBYXKT4QSyJcMLJsynn8QX5aU
4ORivwTr18iO2Jfd6v/UEigLkYFRsGX8XOdWIiAi4OsxXdhfmqSo7FDv2SDb0YIK1Cu1a6wgtP0W
0Yh92D3sZR8uX9oV4I/ajRlo/NCVSaRt+UBzDshzlCnbSZrMjR+nkXUxx192Uxr0J5iPTs1sRZsN
VEdnTzVaSZBGRekmobjIrltGiAp4uZi2mNZ+5u9oY5bnbQw4CeHMkMioxAf1VGMVNC0m0NgC6KS9
MIRXCBcSZeldTt+e3HNJkVuI3n6n+bX6SWxHFKlEhtB4jm05665FDAMzz3BxGQsBjDtjW6t0p4TQ
ODOaAG+/udvj2Tzn5Xw9jOeyBqJBjjoRLJpxtRDGoLSHw3YSLSFaaxfhGiDzNYfOytA+DQGwvn9t
nmfF8LOVV/JJIG+tkQL9lv8puU5OsLQ8AXFh0+Zpc4OuqJ/vWL/FHEmk/4Sqt/jw4mZ2cgiOzV2T
5j/PBkM67ivhXGacB73ZLXS8tQaLin0rKuTk3mJPBQBJlb71mzEOjHLhXm0YHpPjBXYIn7zgB+4r
c7r4qrOn9Zjx66X3RV7FN3A6DQuia+eTPCOfGiuoaMzeppHHNYeIFyU0lRtgws78b0U9Q3seXIBm
0tJY+xUvJnlVmfHvL4vXn9WPEqp99lH6dw3p4YkzP8H5DIgi2gZBts2daNic3VdKWJSLvNKiBXNB
UKidKWw4bWJGnqNjAOhJivRslq4HfhjBzLoiBTnsKMs7P1o1tCiPtTu+rrzD+W22A1yjqDw+iXQ4
JDuK2G0tDgBJoyT0mNa2STfqdyKBt6LqRBngoYAP3JTxmvRmkuA0RrsEO07P+YX4qh3JW8Oj3Bwv
FjTK1qIGjcD3mqwS+XePAe2PqHPwJXks7zXC2fhSrkd2Ix1ppr5nsyPAp0Mo6sJTbsX/cXzE3C86
jZQSCCFZfbzDWtnSzwJoyXHAqVMPYbTlNOuPb96wGxCCCC5fY1FwT7Y6W4ryc3WF9dwd1hk1t4GH
nepLfwJ4j9R2HrWQx27he0Z27dFP12FOfYw88NbCcpFmNZX5QD6nXXR3D3obFm6S6t63TIDdhhct
JsgeNYP7AvmN7kmnmom0ak/KtEklhwo1n1ukB73d9Fbfp2bpORUA8mwCE0bKBwsE0dblxTIbgIiA
Ym67yf7wH0eHKEhR3w7jEHVar9Q/0cE6gKE38Y74wCcsbn7jUFh+M41VAwz4DUGsGBaP/usLGAq0
uSApfSU9rC49byAre0Bnn3bVzvi+fUTIlmeTNIAmJdpaVtOel8AdTVWbqtQw6t/XjnK19KJAhpnQ
gJfd6ZaLODXUCxoUGeqxtvwe8hijyhUyD3U3v8gzBWaoB/4rfRFLbkA8kRLjYcRmywPzWarjC1Pe
98z0SkqBoPlgpfjROFX5K+UYBPwhHK1Alx9Acu5rRkVcf/vj8MEu5AH/+M0yx6Y6eryUMnFcI8ls
OahO7SsTWMOqlbt+GO+AH0Ary7eGmROweUL3tGFYbGeY+Fp8X9lrom+GmmgKpJw/PQfkEQGBKFSC
foaSIe95IYrRCpdkmrvbkUqKeL7cYrCSXxneKjWL8l8CU+GMw1aPvy1hmsUsWk6MWQBdIgSKNQoQ
5is3fxHeWRLD+rUNEk6EGuuyVJ17Psj1LZFeqnwuUv+fakPPXEy8lECHipSd8YMhbO4N+NtOluwj
UuQMT6nziL3lqd4bHviWFe/XaqLOMDGUbWoarmOmkMU7osN1+xkWd/shSkS/w0QgseuqZ5LsIRwH
RjR7XvdaQ/j2d7VDEeDpMfldkzC1SxHjI0DdezFyRYC0XhUgPyhTs+EE82G1yxwc0y7PkbUyOKJU
sy+uYuK7RW6aQ7MZswXJjVzF2srx8NqPPJ02Km8YT8+RFMZYhlwzDUOHmJ/BJCsHErE+B8plfitn
TqxKP0W5prsIVcXpmWYzvRPhaQ0ppa6GNgBHlPUo9QRh71YodXZVfhfeHkKSJmy6rK6nWmhIgTLk
SuPxtjTVE+bQTH3hcIcJgnoMamff8fBO5QD7k1AFsY/5Ld0y9rHQ2asYnZTRYr2CHikepEXxdVLV
L5/aO9ANAHYxyozAdD5QVPbtWXgL1+vq+K1EkC7UQhA7xZ/bWniX7VQYWZPUTk6keEsZWRDVScgV
XUsAW46oCXGT7n4XOiy/IlyYDtZD25yPU4K9nU6PCF2WnX9Spi5q9vqV/SPshDzse/suiRzW+Vgs
K3yHGezxouYKqHDEffDg0uYb8eSzCsyu9A3Z1grTANDNHL1+bjkxn/bicDQr6oXVf3IvkuXplahR
V0DfLKQwVYdrZvZBkBaeEhmG61vlHCVG/0uvfX66k8HNgE7U/ypE5X95q7ffNESUYaQHQFSmSdl8
/WY5HbNUm6RCoty195gTh/HE6dZ6IFNpZwf38UyTnywYDwV3qr3aiZMbre4Z9tA7A99S9R8Mre8Z
/KqgkaMRGyG2I00RoWmExP/KwhOH7z3NVJUrHgyXcMDZoC7HNBFxkJRjEfD/mGkUKVXfGRb1l2Wd
be8PESWolHV6Ia1DqWwYSfwp1zedc7MNARwGxVlgXYq3o9xhY33rZio/NJoIeT/BbM+AU2wcth7s
juz0erLYMqmZa7ADqlmSCYwUUl8wWAUgtbM4RuRlQNpxxfXOLE9kEM68fMDd2msIWJ5hAsBtJTgw
R2sW2k1K53zqpkDKuVRKkJ7CsCCLJArUsHybzCdnGch8XSkwxOpO4qgyBnUDvPVB9WTeZBvLIG7J
RroLc6yg0c4RT1nkrmJ1wXAPxxmNS+9Gh9YQpTL8gAuLRjY+keJz6wd03MJ4n6BDgMf5bt19jwJi
Kw4Rmn8kLNuaW9UMLwb8Nrao5Xzmhqk7vHuXFjRtDODI+HTLzfUR1jLvQAL+ZdRh08Tr1IoYrwsz
UsWPUS3f7fcsbBVurV4Wa3n+OvMMNEjiFsyHtVYMrS6G1dm/bCSqxG2F882oF2k9zHNkzh3h876R
ZKkp6gnhOvKzOoMF98ZqWQ4vGgTIejYgCVk82rnrj0ZbFs/O8B2mTkI3a6md2BiDhu1qRxJC2u15
Uqs27Wt9/fOYjNAY8CuuvXAnS+C8WPspec6bnmJLLaj/+q9TMoiXi9lXOp5EhMAvsRr3JdecmX5j
JPSwANXtWpGUXX9s4Vy66UqIx4r7rr5PGYn3iuajEx+HpTeBY6w//riY8Hl9X/DvFde+mdlZpCUs
xv5u1xkhetDn6R6Y9GNk5dBXCK/UtPomvWSRfB86zCDtB53QcbnjGOVeujwu/sFDR5w6Is9A5MnG
p0BCWgQE8G8SHH9qXDanDXYtt8GtcH2zxEE/lmDehBifv57a+P95xamY1xnPKBDont3vnAFWgals
FkRxPib5n3Au518CMTJfQYkWvACXL2mzC0qNWZGyVFUXMGEP8sD3guE2nKR5yhrgbb6KDFVA4aDz
gtnQAOR5ct8SIzHkanYq/0A56Eq3PX4NoDP9cKntUuKapYrucK0PgR2H2qKGFo6Ab3JEitjSUDJ1
bHPWdZ41zi0LAC224fgQpRgc2YE25Vck2bi41GqgCRN7mFBvxaRI8NR+POv0hK4ogOY4EckmTMf2
uOy598BxxrtE5kgJJxd+bSqlT5OkeANJ0ZCa11J9QSp34+N4W0U9ztrzRVBWQU6m/EtDA+TziNtc
6KkHkzIiELSLFWXy7FsL271544xCoMQLdaZw2XUbQvT/Y2zzp5bMQbMXcupNlD9Umxp1PcnJqjrJ
A7pJbP3SidmWa5cj5R6SqwJOfzV3uyGwKyjKvDDzzDiDabmHKYWtaUNjVvDEb2O9OyTvrbHG3ewU
HHMPppDk2MQmreikIQrymxWzXtujJCQIG3aTzJzBp8rXxtPdEkyKoI8jBZ+RWqvSnzzenknv3Oqb
3O37oq/S+Cpi6e2yHigHItrkE3vmyfJy+1NqGpiuaBVD3NB0luobeZwC8s92NLjAlB61hkGQQm0O
Crx3a2oX4GWKRvB9ll3fHGwsXN90VgQiLDvtTQA8Rw+KzF5YQAV2LiXld46i7OHyc+eUJNtXX0ud
S5sr7n4BNFxorfdrkrPaAULjURYKYDLpZhkFRrSlDjB5Sb2V4GgROb8E9h72NZCydtwTlDA2BNRD
e13YKCyuEhF4SuZ3nhOPc/xwbjr3Wvv0RDgo1zyBtyj3MgEEulb4VxRgmbbdwSwd4ryi5m/ixXAU
YNMkCLq6a3d+yoisTUmXtnMUXMpxBUwEXaaFL8VKJdBYnLcfMKkXBKHCgvmnoQFXaZTK+WBHp0l6
LHC6f456kmrH7pg20fc9QQVkAADlDpc8iSuM8r+3i+z+G5R3vVOA90XVr52S266n3iRZ7Nooc68J
r0U8qn29l8McRZbFnEVfINHhugdw8K1fKvpoWCyg+EkX5WjBIBjffRR16knKumRWzVNrf5toaqvJ
aZq97FR49L57wQmHg6Gr5SyjHxrkZsPGKpCrtuymMfPQGCe9BB4aURGQRdB0E2Mz7BDbhIa4IPVb
TwfE8wEL6vqD+X0dSOk/jCZKZ7OEhvJeKxCgwDp2nlnUXeZeQPyQa4TlBYsH3OoU5gFvWpI2YrwB
+7GS34wRwBCmVd0otVio73d2rn10yg6uHHNm1UJTM/Q42jWbdCfiNE8oK5wq84kERb9BRTZcDZ/K
l5KTNqykQabC0mt93NBSSBv8Rlmc9tvheANV6vBL/4GlAg4u9wh+nKZGjxQXneagorf3+CE7MQ1+
WtkYKITj+dmrkh4F9eY1T7qiRKAOnQGHemp5aFFA3CbF6i0WQcUvTGyor6M714la+lwAPuwBnlCK
SfnFp6Pzv/Cx2Dg3HigUY0gh1t8pzvzVQwkkVGK4s1JbttgH2kjox9FkMFwkWsesK/1ZTdkekCT4
P5WwVyVYMzXg/ufx/zjyDlBkcVZf8uRsptTwXUaJ6lilpWMbzynSt6lxA00Vh2OTbvQTIf9AIZIN
eDD111eoBzb9Vd4HO1k1ZOmW7M7pOolxtS5wLyC4fdH7ucU6YDbEdViDz+5muuNFqXAztpxPFLjS
YxzFrlILIvkjPqfAHBxD83o8mYI6ZgLBaNpUUnRtnxqpYqMd7lqOuK0Wu0tG5KLf+TJjvyFES9tP
ddJKICSMD3pcUu+5yBdZoA3S6Jju2Y3bsMK9qtbbJH1ZShGHr/0+QA0OWWNQhnL/Mh6u3bc+voCx
bu9iZd7u7VfutXje+ACS7z/08O5ovG9tTAC7cYq44kdVfOLtlh3/w5tfOJDx4+kUIabLYtInMUNR
BRabJGNAK2nf6DR0Pe5BnCAkepJIU+MFD4k+OlqBj8M/meIDHYxoy03ssfHj1FUq3pHL2N2a67MD
z8Mth/LO3o1gJ7arHPYWqBr2Tc7LmFq67PGxBNsJ1gFvA6NLX2qW2/unsIoqu8GmS7P8jYuTRU9U
fpa0ISFhJL4XEks+znSi8udZKqmK4rFMreqKz1MqcjY4hac1Bub8eN9SAArrptthP7yrUahjZr7w
AKw/FSnV5GGBUI2DhC2Muvhl3lzMJgaveddyNVtzCRKgkNz3r32tpEeIN1IWudryVrJ9VJmIjiQc
IQb4NqBxIidnqNw1Z0qCOMEKE3JifUcPDWt2eE2v6+9bZO5piy2ARlI1jI9uWspKkVPk5coplajJ
KHXE6gEjLQQ1D+NEEbghqo6No+R7um0iiNFnqRaUMcElyfHSnuEJo12atXdl4LCIScWcOZbt+1zl
qCbbKaOj23hN3VCoSKqbtvz2QG4WWPsSpBfKRE7AyiwJX91F03sv98WJSoLx8LPC2we+zt/ggjdD
6EuqCTFuEHsEy0ybpIGA87gy/FFTstIROmcL+umXaE0aP5JXwcEyJvBFeN/If0ITiuP1C6VeIEeh
IYA1uQv6xXsTe+fe+pdrB4VIvpSFhN1lhRu7h6wwqJR3f/KYN4m8LpmSXogDWBigkGQXJz6Qe7ym
RNJhzMM8pYZUgOIjE6M0cAURvaNoA5L01RujqHlkf5FS3WOhdobe040q994iv2AHwLHdNYGojmja
9azxd3ny0HFZwjqDzfoWFM9Y9CoEH6O63F1ICY2zXw1fAlzFof3iukHIRNxk6BCMu2ehEP1FnTsB
zVIfo6k3YBfwe3+lKhFQVTGwiVFmsrUPeciYThFaMRow9IFc5Whez8/AFGb2ja+56Td0727xUKn8
DQx9U1xfYPnBBGdjNtqTEw5cL9ZgxO0j452GJvTguHQpotgV5Umuyf+nSd2MM/Pb7a14dSHDatIa
zVlIWORDKw2P5cALKbmWkqmFBFudFV+ewzQaYKNnsedhHMec1rDFUWdwaQfSAcqV8FQXKknEhu+5
FxmRDzxLim6eWPlOIC2tNJJAWO/UYT1ooduusks30nKGJ/xdPpbGuh/m1wC4I6N0SviCN3j0y2Wx
IWI3IIscIT2KWqBPkGKesj9nz1S6R6iXJqchGp/h+Ewu9zDejSjAVELbCxCBWc4VUSLIda14hDhl
i3cUecBUaFnoOKpqPWhJk5vmdC1r9aId3K3iMThCCcz5rxYl2GYWtT7NuOEKcPVZbj7laoUnTyo/
MlGMQ86KNscT5ZkXkSD8L8OAExvlcNFkqZelOC1RuN41XXwSE/oQanmErYUeJztazolQXNHkZKY5
yVg04QcbhYvAmO8ySDT8pA2PgJl2WBrGgV12Z8Cs+kae3+dhJzRagBG84zFyjjj0bifnhEcd8ale
LkbcAElZfk1hjCI0X6pn95QG2kJ7hzTNvcBccsTgmjFwe2xa25nH62kbKSB3yEhnpO+pj3qaReuj
ZZt22xiqjvICf3iIT4eOAy/6dUj6je+w56NvKfnO1pAuUE/6TDrF3icEFdqeDE0IF2si9zJfTJpT
4sd/JjHDW9ekVlTsT3bzFLfqRhFHeM0/dkCMTg3ZhHeLjc74gqlDm4j71wtQVmYEbLl9SrJG2uVw
IiakYog6B4+KLWJfhWq+5zDvVTxAhfp4S2lLv0SUlWkSYuUh30JLm9yLtcBgYpoYN3KLQjUw7btr
G9NdXUs88yuYjUVcrraQNOZjqcRQ5eJ4t1pbKeixNDCA4q408DjLaUf+aVuLKFFz1KCQtUQ0UWTN
IE0aSdIFoL/TPtxFMZTqQ5mBTw2eEAukwktHsjlXhoudqizdiaCB6yTAgAcMA58W8VoMV/2tcL5D
PLXqSWqnifw3bs+blHt0OktxTc+rMN0O5zSfvH/E5fvbnq3cK4K5rAaqSH5uB0P4eQJgjIU/4LvT
/XQnJJykKnrpuuTsS69/g0IaVcFrjpfRuEc4i/6Lbu1iR3TK0+uEDdr72E1UVdQ3iZti3Rhxt3/F
xaAIoaAs5sohJ95DcYFfgBWD2ZtykYedquLAXfkR7XSRtKCZ5zMo8Ej0xmkMbrWpVN0nrX84B3dF
XQ1zZiCv8tPOombtYlZyRUjkFdKINjkI0TzicO5fNsDCCwOLpaoeZgfGVt3XrI4lmuADiP3eQ9v4
OBS1Q86BjW4bNOs6EwN24oSXoomuGWReXwK/UZY0Rh35oycE5Y/Jv2h/X4q0BThzIwK5tV1bQkk/
OLmVg3OLAywStSK67lpv5fE8ZTWaNdOYD47CkxNggxnh9ZUTNxBY2fwJasaW9bGo+DKAumCQ+s8y
Kz2rvDpu7g+55jP5kr6IxZF7v6hcq4bXhbJPND40ES20/oL5sFAr6EzhvRraBGSPL600tcFkEq1v
X/sVgMG2EPrmJBL2Q37aqZUp/4omphlh+uSc1r9VWe3popoO/cwivoogGke1o5xRSv3zgm8Yk3rl
jXFFlhIkpoeIz/LjpdHAXJIh+CFg3XX1tg+9PmPuPef9pVcsHT2JUarn/c5YzmutU3rFxJDHaSUf
t8+K9yy1b+vPZIf54Ac9Qiw1n/kaOX8l1nuMDesxGGSangcpEtiy21gC6+kdGoG437TdW1qzYugg
ScPRHvXr7TpxLkjJQI/XxpBANudRWCsc/lT/NG2KoesLIwZO2XOUQABQOa/RIF6UFVbgGjjLtHQ3
m7l/JAq+jYXQOc6T5OBTe55h4wOnTbDs9iuRvR1VS/+VHbM6OsSxyFATXcBcdJ6Nhc0r9vI2IrwP
r6GyCsy6h1joni5o5ZWWTFq7cSgaDIcbhvJyfdb4er3oyMWTT6u7GFfkwZpc870ROQF4loE/N+e0
hvtYRqrN/ayW/eslov9fvi785v3KVYSRyWPE6H+RgU8xeKED5TGML4BjCifE6F3sMfE/2yw32B5y
7jPSMYNm+/Ya8lhtzX0KwP4mwMhO1cLgkHLOG4dN0sBdKlqib8PJxNDjbPgs9UAkvNL8OIGeW20y
4SUPI0YFYJY5sfxmCTeGlRqAqejn+sEMxfInz3XMi5lyX+72FEkNNzA4cy009fbPhsP7CKVw7Ayk
1O7bxLzlS2pDWVn6Qqj+ih8IX/ks8htjMbuikPVZgDRcQJUV2osWS57g2kOZaqCp6w2Ykx21+zCm
BmLDeJ+2QETJ6Poh8m/bkpvWj1NOQ1pDQJHr90Bcvue55n2TgjCSZcWmDNkQHxkZHn5B1bC+SN9T
CU6loQOsYfBuFN7SH/kJPvIRfl25vOwUiFJ1MGgVGnrHCAuAUhJgV4ozLoNrbd0mF4STzd9LfEcf
HCGCs5Y6K9T1MwOfCPBjtmWC09zbO92Ynwi8rXEuJV1e41dYmCSooTdXREhtSFs1PPOFALqbTVqd
NmLyrHns1hsTrgfVKmqHYxe3B0wW7wSSh9l4ppgYEIxsLtix0tY6OZANYpFS+JWd0hNLMt8zj2Q2
hFvkcBKG/5pgzPIpkHZvDwPE1B5yPoJyNgRRIGjS7M8zNWxnnY+yh19VbVcRp33ZkNMtkaOk9NY+
Hif3p/4q1vhbeMjzzpE+lmSqcTi0Ij+th4w1t2RhNNyZjNUw+6mLi0jcyr3h66RioIgiUG9UUNZB
oopfHRV7Kd80Lihs6pgRPClXuM5m0d6vZuIW0kwfbjNj2oCaiAD2oxjzt7ys5RYgNPPyHwJ9Suof
//Xve/Yl64ORpZ/SHtSfKh6Wg+dKennIZ46zA3hZVb+Zg8SdQ8BiCFDLaD1lfyMzIhV54fDFmw5n
MqDnOMxreqdv4h81LFW/uFUs0aLNL6YovXXLWFZbqNFOuiptbtdT71/y6i/DaSi7RXWNg/cDxVNH
HV8m87kIO0y8sTEdHMkSpmFNRvIZYjNuKe3QLNy2aANLNtHk4tJIvp0cM2pRTtPjWBwIQvHzBmJO
t2FK0ffitbL4iSw1uli//akK1Pwajy5zgLVkrH0qI6LM76iVhVzjNWU9GIZwA98h8B4Ikqa83AHR
H173IXrH4jz8HFuxpkbjwK2b5dGL3ccz1dhzS5IhqWopTGeBifOxGzcaLqyYWuqnW0PA8ShzkGMv
m19l0ZNsOIR7VdamN8AfJJyjRY8Vn4+txmBIX+nuKDpIb7x3ZfDZZFIHMIRJJ0x3+U8t3VhU0SoR
HvxP/2zv2ZYy+ePUsVLUVKP7uYqXUY0KQIov/1xdYiAIKBVmxA754TR0HtWFy7WH8f7h3o+2rSw+
Y2upV+0OOXcqvwFCBePz6x+8u9mPzscSre7o/koxmp4J/giyG5Hg8GwQcgAh+5LdVT66/ehORXA8
0H5MlNLID54gTw+m4P2NLUKeHCKs+4I0yYDrWgBXRB7UqR1aiPDdbhnX8K5EcuFSFNmWjpUYvCxI
hKYL5JjRfT1l3Pb/m+2YDJqLB/vGxvOaeoMSD4lskqRI2M9k0el1ZOJjc3KuLzhYKHOG3xqtQt/x
i5PAe/EvzCW5oyfrK0FhDneksWjoLXXVsgKVJyL5f1AbMxSkqN+cE2J1EHH2LwFACAV38XouWloJ
x2VAGD89cZhYcZlZda+uyuk1mXdYOP33WdthptSBXRsb73vwTMziPwVe887cpo3CnsSOnocx7QQb
p2AWRbAlQYl9GJWTQsLbSyLurvtuZjb0YOIZA1MB8ve2YAZwss6u6A8vtshKWHdX0KQKbLeQyeV5
ZE57n6wFyvgq2sGEhnRSGo5yMv/Lyfham/qzzYb8gYWwZHBQDpuaxajz45hbB715ua4XYjE6fvcd
mN1rxPDKeITp5x0rc5Or3Aku/7ErNwzJL/d7A7qOUsqwfM0NeA7Hg/cqvgQRZ9kmyP1sF7a4mm2m
r1d6he8USdUovc9S0NH6r/ZHYamw1OWlpwE8xc224k0mtCmcXGE3o78SKEbUuCOSmzoC57dDxFv/
xQpK7CSnKmI0/CI4ve8wasTBOfhOjZQxcFRsAiqaOZoE4f2l9j65cEsTS/pA2oSOKUMHIUxcm+Gy
cmF9YE2r34B/OfNSSyOS0ql8ltsJqaghSBJpTVatVHFwvRGhZxuZUW/LtOuHAjV0f278YKYULd1Z
R+Nm77L5vmLTlUekLoC+HVwElYO/FB+pXL5ifARwZvQBaU7HV7NOEmzZwQLBKRaSjPjEaiJXoQgI
1jy3eWU64a+J+5lD6uBYZ3JxFJqLqF0RJW6GITPbiyBE4bCJIwdiwH5BEUKjwviiV16z2Ttd/vVN
OfPIhsTLOoYo8t4SpC05ZOVe5G4yifpZT8VhXSNW97oTyPor523RxavDIU1w99qHQv/uskjvTR7P
VeFCQoXPL+SVxAEu4f40wC9PzP6Ge65Z8my+8WYBKmEqDDbuPFxxpqPxu7IyIdnrJYFw27v5hgh/
ZqR5XrvN6vBAI6uMuqTU8EH8y3wnV1N6u7Z2kxOC6jHtcGgPC8ELH0yTgda2itLCGxWuKSJUxat0
OGpzaiGee9r3whtp414B7qIw1qRveLDUf1Dlhq4P9J3aseyd3Is2fI13m5RfdlbH79h89oiQ19yP
69jV6DKibnEQlAcYL5OCIQ2lhjaJ/6P9HWq+5HhN4xAuwIipcVkzjwwnJODBkM9z65uWZh05aexN
BTrWi29AQO1CTLlJJ8chCrWC+FWGHJR8p9aGFAF02FzOMsnO7P5Vs9nVLhZ8xcjZfD2+w2E0M1aa
esibaBlKpeaLdrvEqEzmZhpAVvEpj+2kD82SxXe95HTWxMls3H4RmZJBpJXrkMGFFJGjM85z1xG/
4Y3J17+yuGpee2mLkclkdpocu0OiVP306bBi5/ZARXxX24eOt8u/zgjhhbJCp9Y7XzyBnOWV9qVK
u/SfxjTlNtZ7rR132hYwfuvytLaau3Aj9kyMP3Id7ifOaRnaJ53PlwSh2bMS+Qw2GFSMejWphML4
GPttX3a2zyo98R0nF25zSQ2WDeQ+DQCs9UKzClhc1ISOStE0kKl5YVqwcIU65cGVDHtxPzIJNFX0
qnt6eOyi70W5jpVlVhuP0ce/lDkJzPAnwlvqvhgVeFbz/r0dE6K19L610bMw6O5SyDOQuguC5sea
Lq94IEmchlnTX3eSLx//t2PFUNein5zig1/++qXeIp/8Oq1KEREImCmEQEP4ECWSya2JBYvTX8JY
mpJ9OYsWZoqQFuhStDKA4xE5JeN1C4Ikd8f46d8RE0BwJ/WYZN7dHHxSdZ3pEbliTbXM6E02QKLC
g/zARpLUZp9f6OKsQ9klIz2tCK1MR2riSzWUOVUt8fIImZkgg3jbyU/JVcgmCUpjeHFVbWrQg+U0
Ii6mWU5TANV90iutfk61EqD/q7iBSvXysggexCUOAfYwKADZUU4RpyG7UoPVqhxeMo819loJEfSe
wlQe3SDvAOZvF97nTI93/hgMaT/2bwDBqf2wO97wchmRq47zCGGT96Y+ZPdZT06xrHuaeLP0iEwz
C+b8Oecr0Q3trRUqQZbodZloy892mQimpZdhRyJQdVtIIaBthR16iOitKp9dwFXu4Knw8pPS7Fa8
icVe4RbM5jkHfpyQw2zLDeuoSH2Ldlb2sHbvBM9pjBLsyNHc/CSfH+m2yzsXz8eTu2BvYkMWJF/l
ukCsCZDY13/7k7CGy6sMOPiGky7Jt7LJdeCWK2WiUm/KFTab0U2rocyg5/aKZxUjYWyYVvnvJmBJ
kd3w442/msZqbiQUz/dD3eo3D2y3Dc6+HiN9za8bcljFmRSaBQN5rcvz2HceNtT2U7JqsJ20SEP/
3rOOQXl8gf1Jp2GuOTg0wQXOEJVADAUusP1l0MXrImWXtLi+o9MP3HDHCSZSt0ZxVkzn0GNMesrq
qCizeiHjVxEP2lJ2fJ2aMcEgcLS0M6oNzmnMntxUHb2ZXgSGDu315RJMOdJJoHqfT9ff76M1m5e6
D/SS8qaeppSz0gHlHypPKkSVB59IcDMm2sAjh2sw9PNInosVRBLaCUj/UTJ74QaSzpx/3npASaEN
VQVFWnf5/bITK7bsyx0cqPVLtFBBmMHUfWSsNjxE6aA0zD9bRob+XFanOyoZAkT3NYMQOe3IaHBk
VnjVU2jG+qK0+evy86jXU1q3vq6ZvyCOpMtKfv9KHjtaOs3UZMGl6J/s0Hsp8Xfcieuz26bOyUev
Y8yieFRHn8vY9yVLrILcJOrT0POnYwLv58StivQSj23M34P4pAxZF4fIf6P5C9IRbBtXGhecD2cB
2xz8GoWUneFAC2f5BOs9+jxfO0kYzFj3yU8Vt1cNTLpsHOoWgkUfO/+Mw4jLMM0PS2CL1kjL2nne
QlAhajl9jAsSWplOo3UzasuMe5OBw+ELdsoaRIsYPpKe553qCzBtx4FB8bKdhvYdKYt9mSLZydxg
zTf2fNCl3ZMXVuuIUkV+a7XwyH8S0wPwt3WUnuW0m5bpg/8e8mBB2HGHVVdG0tA552GRXVw47XxF
RIESOOPccdXkeJTIaeXkb6JIlnwAbBpoOnqLONY6UaYJrWTMePapR/OO3wfTwq0CwVXVH7UXKzBq
X+BODmz8IW3GPtUZvcWCF+b8wT0QNgfXIzvG3uJyfglGb1Aq9qG2F6Uh9b+ojjgK9ITZZ2UJAMeU
1EguPJautW9Bx0O4J1FR7CTr5qfLNsuwG3DEpTvHXzBunTDogE2F299qmo+b4fUlT/7ZPl14jjPE
Jivu96R2q/WZbM+QvlhgF3pr43cMKSbCLvaYY45DMo9MRqsof0c+QQZKJmSRBCvAL3v3plJTb5JL
XcR5Hl0NgcDLFCB6bbH6i+tu1Zdsmz0gioDkhxsK7ekQsh4AMnRFcxsln3JGtg+4Lpgls55rmjeV
yv3cYc1KddUxuKMz1h+OIGdGKOLAkJryJlaN/QvewhlSvLzOcd5RdvDCnM059+Hs7pHONLQZIezY
jL8scSPbJyFfj7fD5s3SeeC3gIsrnqMtY+bLGZZnrylQ/KgHZW2xL22DOwInZ0GX8KavQnt7MKYq
Xtkx6qtCmulV7j/omCKLxEh7adUpOAFLug2vaOD6puYZQcEjqnM8NHv/ZcY6Fh7gKEE3Bbx/zVTz
Ugm7Rx/U5s5Osdw4PzeBym30+UpopHn7QvAN9CsBvv2cR1uZRN1q17/rI8pXOiBxG+X1TACS3Xnn
NoeWofOaxHsuLiPdr2cYgdHFgDoo3jpjoQ3rCbhWrMun7mhaJALlDVuUMOfUmwa78av1tgLF3Cek
1uhfMupCBAXDsg17wL57E3+pAYROYGlMDKzbm3Nom5ajpFvrXXbWCa2WrdXno1oHVsLG0Rj+Qrmr
RYQKBPktZXXwrR5F+7N7Zx+ZO0bRy+glk1tbDmDjpZVUDSLlkZEgkT9nqW8VZW01lfXZxYF6xXz1
8xbstz5Og5G2g6eFgImrQ7WqEztaOn03fGX2EOZnFkQc+s7HUQmcAuZPoqvIExYtfJT7WWqsCrmm
tT5x/vCchLkueWpxYBE0ranymuzEtk9m0s+y5b1aO8JCFX9v4oMN/LrBsdNNUPZE4CCayeFp5Jrf
67zBI7/+tbIqjbCmN72xBtB4v3459D1YhFf0FquvjK+mBlP1fLXbObwq411egsfpyDNGh+rN/It+
4X5CemiHK7TmidbQZTNcmB/0J2A/WgaqonkV1NGCElgVGihti+Vg/J27y3VNLgYaHWkQ/065Ap3+
QBfas2lXTqI8TnSNKncpsGFv/fC6s9LYSwRGPGHxlxLVpiyAOgy1wXZX+MQdIprdQzYXqGH7b4WW
DOPwjLhvrcgxwqVsV5qnMrq+BpUPbAxwTUyDK8QWglh2TP/1CPNsja6KFHib8aOl58gR4Ttab26A
zi/BEm+MVV06hUEneJ2WMGltL5x4PUNzUcG4YICQ6o6r01olfP9It2QaG3YdWXl34JfB9LJt1rXl
PBfMhPzgPo5Uq/ahdvPR6Skkb69Gl5Z6H7FHsXfTmf1mmO0jQrB3rlbNo9nl2jpJpccjOHKT58T9
31w8+oA5eShobMWi220ehlpEd0k/ycDhZhhs2j6QXHbZeyP0dUlpTPevfcIEZn0eIi2QTYiodosT
FXKkDIZo0R1yMvrQ5iZwj+IXcdG0TkKxHbSo6SeYRMsETYzOABmqL4Hk0zhfAtWk6F2K2VsyRU6X
ymsL2E3/2J/EwW7lCODE8gC+Znd4eoKXHgkj2xwNwtv3VNfz2rul+x7QpxmswHiI+edzqxjE2oMg
ieVEZxb/pmDmMjN/V06s0gZ5/qhRKKYn4PM0Sseu79oZ3Grce0SDJYihYhmCRTmbImcI0E2C+faF
7DyLg6p+TFmzscslZN3LnB7ivL7PljADroMOijliELuFgFfaqgxnKyr9BDMEAVKw+9sZ/Eu1vpTp
pIMz9mVb4rGNJN4J1WPtZqsm/DSSCE5yH+8oSxHLmAgy0lvrGbhmRhfJaVfF2WvhvF+QBabuPiNJ
PlkXsEi6kAUJz30OZmOj/tnsl59hR5ZqtJnd2/8vieqYlqkg3n1PdxJtcyHQCfVNcBx1y974w7Gk
wjSd7XvfkJfIuBhIA8WzRxNv8xuywzFHxApGW9zMTInlVw7TrEKi7qr58vMDfAYCzbDWxDaP/6WN
VaMuREgrDGnh9gigaqaOUILz44Lh4sWmAH2KBi06sDnjmx1mafKNxTCfVvqYzKUHcqzRKhcfFxHf
VHs96fYZSYgV6rYbA50Z8VUzMLjA6hiUvkbJv+5j65TSnuZu3Z/451wIwPxdQ6+5Dx8goe+L9+iP
XKFhgOx0N7UT9ZoO0LD1jIg2zZ6/dmqbkCCRfpRY0IWQMT53gfj3JmKik23PS3cYoIeD+eWgct4I
YprGuP0DiXryqOgArqIAxtERgYGhINkm3Wr2sQlED6KcKU29ik8NQqqzvOCIGcpBIu3CvB5dskyC
wlaMbxFwEeHYOav89YZfxuvrdVFsx4pd0aavBgAyHXIDVFRwJeNjq7lQD1WKw0ylDF8mcTVX2HZL
K9Dlffyj/qsDWfNRisDVf4DrO1TIxW3jM8Xts+fHMQufYZa5dF5eckZNJZQ5weYq1ceBB3RDN5+K
Zhtm3NWBO6ptHr7Ti2frf2u3zxEJdX+MsgTPBhOu8u1Y2jY38duRcQvK3JO+pwOfu7Kah1WEPcfo
W9jmNqz6zBSd9zPr9yuqCb3pmAcXdcRmhNfzKYZfuoXJrdwDI0Q/h+ii5HlSFZKPib1q5+qVPW1/
H8/z3zmsV8w3z1905Y9hasYp1wf3JMpvaGtozi3VPdryNEeaD9IQHmm3UXDK7GN2d2tTpHRx7MQh
Y9jpQCb3hpTh4BY6tPpUYJKvSY+OP54W7ixyvgK1xOARCovqQwwyivoMudMhpC224wo9x4GscOCf
KckzmFCK2A9D+9/4xEhsv1vBoz10Bu294a4OBopCwUP24j70CLJMSF50+tO0bMzAdqJngmLmY3yu
Nr+1Wx6/xG9Xu4PWwTYZ0WrRnmFQbwa0W4JBqVzKX1YJOLLqdotmTbmSOVQwauLI7MJKTf9d0S0H
J0dS6qBNWptReJme/xg2j5MqrfL3yrOnEX1y4jKBISIKeikK4JHZtOmIr6xxDTKhnO5LpRDR1iUZ
rHtnmnCjR/oXzgAhFvJlkISRP6krXlA8GgHg9QOEPU8BrIKkls9wrNA/PSK2B1ox5EuEGx8k8/VN
MUo7Hho5USUvxFRLDo1k/ZRxjJn6UwWxJbtLC17WKMSKFNpYTtDPKVVZWaUJtHyQeQ/+qt+i+VdP
jzKTUJJY9Z317zmRhRiDgcX2qc77xTKEQBg/3eI+lvbs5bHaLL369j1iPhtM6gJDQWy6cOHKywM8
CMEx2DXzGQ7GnupopAMxVO7kwJ26EhQQgnDivciDiLzLKpBrDC/mZ8vfj1rJ+Xy1JbwcEenNpx/6
P1So5eHFmcCSa/W1+6sJMg9BP1DMKpD+TXf76ZSQ+T9CWBgYF30zpxBjEvzNuAufIUK5dtnVGOv3
2hFEaHTswnvl46HmSNzE2aAmvWW94XJv9tQBA36iE5F0FfwMbyZ6H+6WHDcakPQoJK37WUEnutIv
b/SZRlOWHA0CNVYmWq0QW7SDusvW/VFpFabgCsPYu6evAZSNSDS85WBCXBZSw5akZpRbGOAvWsYc
h4qsphaH4Z6syYhvA4Z5P2qysNxOPsLpBr5uww6FT7HNpWXjM5sL4mp9nXLcDBuC5BU+ZSsg8kMz
JqPQiZ8dyDUF6U8qA887GJuIVlxGo2yEj4h83d9M+OmEzJRDXaiqEmNyHdn8ivU9MPPu2oiUxZv4
lXzKruQV7GZZEonOxNf6gGlN+htPIn573ZOK8O5XbGJ3/AajUoY6fBXhfRkQz4rhuQKffd1hle77
XnqcA8W26scClSXcNVCLdmS8n7TFWAWpUvo9oMYDiPQplzXFLXMEz7ZyTHNU7gIoiw0+r8fGJAQn
0KR+Mp8I5Q1dBgWXVMiU4Hld1FLcViTHaxi13lFZvaKNYhsnOhjizx8ZbK9aCDVIPT4A0Eypr+6l
dUocYZyFJbqQzm7HqYsZXrTjc3BCJasPq6Tz9Q5l7ZqDFsPJMRMV+N02oxT5ILCREO4SKfC25HtQ
eM7/wgQqf9KB7vXQN0SOfUyWcD12EEdetDYKp4mRypaasdM5myFqC6UpYBG+IuyWPsR9X9EvLkpu
maIpC5EbuqndCASBTWfKIqpV+Q2+YGzk5FNIYoJKEd2EkZ2T/EOWQt6VhN+09ah9c6irG8kYsQM6
3vdUfp34e7N0GQ9AFHcVwxtfHNdm9nZdi/YhLZn2fZt2ovdAHSrjmCSbWNYRPvIYZFaasXAz1+Xs
iDO1XDt09nQcO+K8RLHHtgiSeAsM94JIwkEHxyXTii2+B/6VYPtiVh57/Qsbe7XPyr5L1XYmWeQb
n+CWRzShX3P37bbO/Osx54m640Cr9ZxeEjFG1WkSr3xxSHJJSuqJoCMRimO/TeKsRxj/Vn6WQdla
x7dBNO8G36IgfhyDn0YJTZFk8mKgHy+TJopTIlZT2IA9RB2Pt1z1tLf1B9w0YuCLoPy0lu3vAg/0
fCLUyQ7rQDte1/rAEcIY8cielAfgy3CjhMmoXEwVVQxgkT/YE8FET+uATRfbhJSgFe85PJnJURda
cZiuf44EQem+8+KxTGI+S53ic4gojEPpOx4yk4SkOqB16DmR5/8HIG4Js8lOtNDZLU8YQBgJCS75
dxBeDBFbCiR29IIUfj8s0P7As/mW0J1EZUlsDVa/83Ot8rEnyc7uA2HS7WNPtPUQKdCe1o44MPkU
Fab+WcENfsdPDgNwv4QpYngmAL7PbpGHaRbURRgasNq2lKz5X2Yf6m2AUv+GBexYZy44zq5GBkn2
PDS5MMhuIbvM2///8ff+KUmqIcbXbweOJvEHSQ7tI+vLtWPP8ImuMIJKT/GWDksfzmxW43L0hqxw
ZDkMbp8FeIGd4ySxyBZFGUi/ZJoPg3bxZGfyuH5+qrKJNL98Ks1Hy+wRK2llIIj3kSIuesxJV0EQ
jL1nfD0sKrwYIYbH3eNQHaFMMUhJwqEW7YkmPVkcS0nlRAx8qUcK5yFYhxyplHlqwasx8owBwoGA
SAGKUq9KLmO1ibsYzZuwaNaR0Wo+5+bZp2fqgqheBdObYyHbTmucnQN8u0aX+VvkumXjzjWtDIy8
fJubvINEZn2FK0Lduh8LfAuJTX4wGNDHB741CNP8j3o1HVbruOC2N4JWNkYYo43Wr6ers2hQFaNu
Rbr+l7OjPRIjyzRUt6MRDcabTfXnX5ES/tZcJZLgCCW+YYj0E5XOFgtmsMODuUcjaZSb++KsNDHK
kclOQ6UhgYI0+eCrBXm7Y7kqKCO2lKSay4BYzhlOWi/ZaGUE4RkxPrPg+VyIPwvrlroWAj6VWwu0
grURTJoAxZfBV/httGZ3DzsbDYDEsgjFBn7cqvOtIAjRtjz0O/o7dGeMp6+zUmx9XsA036mbnQF/
4WjCzyeGYlVxiuSZYKndHIM335vWW6CAKPeU5rlZrzaxUMD2xEXs9mqh0XBNxXe/SwCKF5XQvxwp
rX3ADzWvPH9PdoUzNzoP32Y+5170sUBHJzvL6D66DIM9iIhRYGsyizacXnHt1/4nJ+zaAL278zhs
eMkuDEP3oWVABfu4EVsJsbFJz0roenHF3i6sFAly2R/5RunNPkfucG/SLBavRTddgzSPqiixJmeG
iWbu2CKIXEgjCGzdAb2Q631fSiOFVYxtgopwKL8yhAVQIbG/cbhJC87ROk27snrgjN9marFjtDMV
6e98XS1VyqW269/nyE6UnZA6j+QF+dw6Eq3ZKW3N+lPXZ+lQ6tAqsj2MMduQoQ49rTnQgVXfWsjw
C7eNTl3dJzZsTszpV32kWWDIguVi/k6ogX8hmFIzzAkT8gFQv5te9lXgjXYs3J+aR+ryKt+w/914
JS5qqP6UPFP1e2Vg9k/n5L0a/ZM5gk4/dtBUK+qU+DNRmx5hiqX1xVmT8DBRiV7vcmApboo1WyVT
rukIKP8e3vBu5XggWacYOlDioGWUqf13moR/JCqMPl23qy83Vvu+CbSaE/PhjgfcwhJ///nqn2wW
XHA36Dl0KcXaDO4D4znchlUXML3UVTO2pLQjgUsSphNWl+EvwrS+LWfm5wvNtobg2deQGMmxAry9
6CBtZNd54CRjZPVr/BCqdaVC/t2+uzaj+WkDTPM14nhm1If7jiKvU8tglwDCk9JB+Eay060SCON6
czr8y9vftxbQAtLu2swKfqxoYwLpEeQhjg+XXlHoaMVmO+sboGkD/eyl7xUhZNirSOx/8BPmC453
En+K4E041XOTqx+gq49K1UT+MzPxUOsvfTTwhPm0oyBwxF1gfQXfeNq8miHFBTYn1yaU/7/TLaOU
YJdYirBzGmTXO/2mzW9V4BO7qGgox3AbsLjl2UrgFWkn3qXwpVPt/f5+9XoqZFWol+4tV1DuyP+S
ZNXRCcYBZDR5+/AX4/CQykd3pC7LKcFfpIECHWu/pNhDUOwJ3+g7JsstaJko2svFIu0FfxpXNUnj
/18hnGKfFxY7v2fkNpaNHR9xL5eOTwLY79hhUq4wchqd1KE02wE3HFoHG3EscjVT2q8z6sgbRelN
AVjTjYxxNhdEJIA5zi9Nve/pUWwZSv+XdQF0CMxWaM1bbDZnO1PCDc5ySjWtY4W7PUE1BNs5unyP
nv1AlSChDNo/DzaYIxW6D0wkEwC16CwMRQz02dWZrv5X5w6No65LoqVcXzjEq7aX6x9PojUEaCtj
Ki5sF7wGzdjT9CzZyqbXRc4IIW3+G1d4y3HTlk/5mb9beS5SRP9zCXuVcqfsEnGroyN08rNylybY
wapG3OR0wkFYxQy5VqLdu6oyjzKuXzwSVbZtfdARimvWNjTZyrhNJpqDAxhfrZFCE/JWm+aJs3Bt
wBkMNgT8du7uyLlLRN7kaQM9/opRa4sDM2ppQncccmz1U8yPEZxnlGJzhsI+H+2L8DncdgRoPD64
iex+9e62iCXzIGkHkjziVbzwAARW9CbPU8CcZg2ZIw415h6hKeH7Gqbdgo1CHBQfadAcrRWYgJKx
CnDsowDhEdzqRxRuZYtVDMtx6jI7DtoSePuaIAuziiWzDIBcrjTR8eJCKHvUes4j4kaNVGvhBIrX
yY9OJkfXtqOo7epBeX7PWYc3gxOnaYbCf2x8ObVg/ZwbXv2T9pfF87c474EP2k7uGFP6GybNfzAm
Sx3GhfAV2kE0tAH+9KV736PVhQIKu/H8qnuDFh2ylavv9qKfQNSstYf2Nb2dzFJ8gBh4YARqnD4D
4pEg0DyVRhM/7M+3mqBgUXHOjvRVk9FvEEUEo7YIOQ/cQXN1SMDLYVbW3lORS0b0lAHJfJL80uq7
wZkkBihfrgAFGDZHyHUFgiqLteJP63YBgdPUyVK8it5fW1OcKHkWDNYPre+3x4ATGsIEKzH9sXpz
V/pVg11awmqoTziGlNwvcOZYDiWrt8g4ZWr3wJXRFHIZlji29rqqW89t94nUvoRGqpOftZ/k5zwc
ZGLw5BcOgdOCdaQE3nSa7z1m/zEkS2HyK8iSduW/5VH5qY+FhsL6CNjZY1Tt4Y73pFhurDit8KWY
vMfF638+qr4RcLmoRo/v4V3mZ0bI08YAnPqxLpojhMMaxyfrSd4g3DP/e2q9dy5W++0JXqPMkEej
EJZS8c7GAVelN0L6k33o8alvFu49uP/MsYARuQqHt7GNqu1jkkBh7sMJdNjv0+wjUkH4qFLyXbWA
xDpYKaJ5vIG33pToMaD0CLt4ZFI/yBkAQKDc756VD+MZnoSxi2Z157sNhcmDq3Gs2g+U45v9Cg49
23XWpcwc+nlfSFtOZaPRlcbP/3XMjwJ3ErUFgplxkNjHKpBGlwwtUUN+XMJEjiteecClV0tq/zNr
5bQ/x0zpVcRV3ZVrG8AdknByr2Q1IQaYSdLWgKuBvGqyh35mZo7nkpn7oC8PyPQVuiQA4ezsmaIY
Xgxc/OlpwvIydAXY7yq7SUNClOmzhS4FsRsQZ3sx+gTKx9FYozCCZ6ptieE8RHDE1xqXV+w6YP4v
yiLp76IPm31I38oDa1IHUT3YoThrgFLKzV/K9O5ottVUUDm1O10KtPRkjR9aBzz6KVbHkIFGhE5W
pVehGGZWZM2EtlofBt2zxhDGRR9dsT7ZUGqQOLEqArOhBO8y3N+Ykv+krTxHj5ECT87Cgk5S+FIU
GEUJYBge8T1dVSp3k/ZCCVDEHqqeKC7goTPm5qhYYnFeW0tla3pN9KnviqktNW1cn0q/uzbgY6Ib
dzKrUnUIZs/XdRBuiALmQrzHHvCkeBWO7YLwo0BaK3TtgbAdQp4wLseuMF2B1iMn7tNJGQHMge9u
Krrgbr0qFd/0Bhxb8eIlxiNGCzEbub3pALeOBDpe5fbU3QMbf5nb5rUGiwugwRzIzFd9rvIm2JNc
kPNBTo90dWj04NIw1cA/PpyE/ip0HjTSiO8fK0mIYam6vXdx/MWNp0P/6USHJi57TwkzOeGrosYv
5v9gBtHDPXNPkriVXtGFXXr76GfeoZWQxgItIAmxUZ8bP5xjFgbykqCByFQ/wPtYI59gkQUvUsQd
aqYJ1JeAW78536rY4qVqSF+7V7iH3pqK+n+BhWg8qSCCGg8GHsvKQNZ4dwR/S9dqLVZOb4UfchL3
QGVt8LlD4KxaS20r9lVREfO/0ZeGYFtuVC1JahwW7DFxMItS1IbZTl8+YysAQs166J3NWNsAXhHU
4Kgri08J+z2RdRy4jMOHc44d46nX21jnn00BQT51J8OsbMYYvcgq9MDLlrM5IrY11DK6nLXL2BgZ
6f3MCfAeAthrDsmvPFtxufydFgQ7MG7903mDQXxQLf5G5yciSrVRqDRSlfRPQ5oJduyKKtjAO9uI
iuBAASbZ1kKNPBhhl3oM0bGq7wqz5Yn/SK9D3FeAyrpeb/meoGDCj/c1e6viXvqLp6f8L5KcUhvz
HSycY8R8WG0wmK3BcSuZR0MO6JqFd0XBoCDvPRf6oohCnOvCyrevxEOwJUjOGsR0RztL/paT5RF7
2Veor04y3HK3m0oe8832TWCADNpHBsK1dcZ5hOoCaYA68jtTwHYPeQmpB9gA5ZqVdJgWnLkry56F
w7tdBDbDmseNQQ1vPR7eleHEYzx5sH9W09vTNv0b31J6WfRpJ0/BSlQKtmbnRZHflnZD+w9jA7bw
qOZm125sFK5jGgO4fNd9RD1yPTdfp7/58MskVKMqC4IdZ1EjiosIs/XdV+WLkH9NLW+CIrAlNuSV
Ylt7hyuFelTGv8xmE93kGSjkP03ZS//fAhgvAuqa9mfJ0RIFRE1K85MLqekvimqSb1WgHxceEzCq
WLOsA7f7JM5S8lZkBg1U7E+Bhz0xERG6731bg3AQIYJ0EV7yrggK9hKIPiK5j2Q1pFiziaVctCda
xq2gXl4NFaS88/thFb3CyVtWVLFhCPnAFk/8ZswUlMsGL79xYGueUa6AF9YZ1Kw2tXhCz+puqqyH
pevKpKY2ZJQuu8RQSsZgh9CfqVVIYwGUISkn5x7eWXP/KbKIOBNCtUPQJVot0ltLu3b0WYv5gLCE
mfZVUx6eqZncqBOnozw8S4c9aGO8qmIf8kZUfelI73+4djE+L/xaHM27D/OwvJhgPpB1TUTGeTMs
ewMsiCg7Nj58Atc6w5/jae3OYTLvWKR3XuuhjOWWrCCTZImjE9JYQ/JEr/rtiFExgbGBMfnNroAu
wWrWKWZAlCcdE67xY/FD05g6jg/07LPXGvE7CPI/uvJ6CEko/q7bfyp8iWktvCLAmZLTm/jTLprd
e8vQeOV6ven/a6LFGZsrv1rFaGckuBOOgI3Pg3m5RsXowdLNvo610f7crxqRi60oBSXz1t+Rdw0g
hB/0l5ptnFj7FnoSNQOiNTag8PX7M+NKnObWR6ZEF7UNATSbDey5oa0owXfp7Kuc5Lu9tr8CmS56
KCCnzPs/MkHEKmyUXo2HBui/OxNyEXYKYvItdu2mZDhvMElKuqCxdAmh8VYxLaXFnjw9sZmBLDUu
v1vc3WbvCjS76LkrBXcjT2UgF+j9Nn4n+h+aEjd8EID59UP13H78fGuM4+SxOmPAd8S3F0O4ZUix
ZGdOTEFctJy3kVDCyifauxYu47jzJ/hKGmElJ2VIKGiJS6HNcbIxfqSo8McAdodYw9UkwezptE7P
hMNlyLNKbkETwmDH6Axu22Hyy4sG7FRrbTbELmIbHL1zFPm2pLeu/aKws65nYc/2DdPUTtQOmTpA
vrrjX+gCjdMzZSiH/2D/z2cJ30JewPiH5xe0nsVFGZd5bkTaUYztZbcW+DJGZt4xXt9LABM1m8ME
WJxMJHncUSYn6z1MUF9f9lvDNTx5V0ULCXLQrswS+coviyaIXDBzy/RG8dZMoQy0FrKFlngzSCy7
5vxLgy3tAxidRZJJO2Y+YLTBk1qNu1/8wH2lHiry44F4UCHYvNR01GTbOkp6WTGu61f4/F7xG366
3ljrHENp9TjOVEdE6MjE6/SOPvg+OcY7UZbURgIxkOCgbapBW6rV5EY7hBEmY/j556PxvXcrGhP+
jap0aUKS3JE5zHueDqXHA33nLUoFnBWoxpEPuLXcDzQxHE0FwEXyXIibfyi5Ji6mPrnuWUf6j6Lo
TjqmGSd54fvGLonvhsS4a9aWr77YVuoAjQaxyKgVnEB7UthuNUFNhhL7yNjxDAXxxZInJo/PuQ67
FwNN9naJIHINbWrw5na6cW9SFHo1PKApTO55TV5CtdGGPeQRg9igOH5Vz2QbGpdWCNn98X45qLEh
L7F8gf2twFKOl40ukjU93SFg6UHnakEpZTaMkd/9mi/jxGC4cxrCyNRiqAVjqa9cBgVE0m5qlfJh
TOrMeidzHJSI5dfWoAHMaSoYIjwBf9vvOPUosidVN7GdzjTvJdGHF1Na+D4CCtBHsmhfIB8F65/G
XS+A+rSgv5rjGzU6m7F46+piepfV5qPN2iaOgWwbqaY5+3GO0AGsR+HI+akI0dsU5mOEBZ9pFnq2
GxwTbmE6TdjnKAiUO8a/jt3qhBRtj6PNYpgCxX2hdUlmhg2sbJrUyy7TPzKIJBH8vKroe0utEWbL
TkLz9uuGQciWnt1wNXDL4giDNJiIc1Um+CNrI5WlgdXcRDAT9hlWiw8FL+mzb4Xy7x/p+hynBKgp
P4OmWuPF+46rMfPe2cRNmSW1WFNRjWjyjxlCBxw0NWKUM7GBziaO8k9/1VMzqxnn0GUMX+fuYjzW
rgcPv/9whWNMLbqGMMQydf6yydWVqMFwWiP8oss8bG5sUM8bVXz6jZK4w6YshL0lFb8PN7CEqtjZ
H1bbzbrXsx1VKvRYNvqmZ3KUxYf5q9PmdK/lJINWB9kVztzqlkMKKawjWg/n6BbOWoy2xmsz9AlN
tkz+YgpQ2JYCLOpmjGvv72xdvQ5o17RILdVdeNXly9kNyK1ZQFR4I0LCq9FJwIK3rShB+E8hicnl
4JFcugA8uEhUaRcA+6OppNWkeaPdggyYpUIpEkFKQcphrxZxplTvl0hyZegwcZomkqmDlqK+yWlI
WUqzYIxnhlrKtli3IlnWMG2dKkLXApMXY13xj5FDfuH3exabGS6ppiyBWLi+/0+EI/B2B8AkIieC
ZmI8mTfRf45VL9r7Nhc5pkC0XFrsfdT0bqWXWWGDjqL9288zEsPCJL3qsThLu2oePfGAuZfGHjOI
wVWOfOVJ6uxxcg8ZyR8ReVvCqo0nfGbB3qRIDJrXiRM6eErmrm3Kjrq8jDl3fDh8EZcpCI1R45bZ
tNvg7I5UhSXBGy0OSYyeIZNsCPO8JzBT9h0xl5H5HvZpjTr/ngd25uGnk1ZwcyU/AjjT59ZivmgM
lJ7dCa8mvfwDHWfxjUOMjuyQw3Dg6I0eqvRqEpN/hB3OjyR0ttmh65h5UhsjqPgMMUNKGv+J08gn
z8CzDwHa9mEHj6x/SUiVAuuMcV/0xyy+QwQSeOkBIo8WPgyjJ/HGA78YajQcEuAHVT4uAsc+obDa
ez8CnS3fCm77xdCNIXr0q0QhJ0CmLzBCK7t3wQ3uE5uFett4yxGx9IG1ymrQfwo5fITkELykEDqd
vxewIwRyaA+TejTo0JMhI4S67fu77yWpOYH9jybg6qikmNa0Jozv5bx3ctAGsnhu3dXSX19w6YY0
1o/xPZXORFLqmywh2IFmhRmKziVYpRtCoUWre/NMdYUfZ7a3xksEiRCsdbEhCLeHm9PtH52L+1ar
LNhT1amh0T/FnmIvW62TD8TI0qbFMlC0uIgLRJ54z9ySn67ofCJ6uTDqvxSBAo6Z9PQ9bQvWLCbL
IPyP1DmmLrUbC7X67VDR+5rFS2mJnjY9WzdYdGx+Wgo2Wb99L/lKPWkpF/xFIcSPEJkqDFWYisNa
GzaXrTngqAMFPSR6g8Wmpjq4zLCoP7Lq62k4M6XBsU2ZKmJOJG2vkE53yd0KTJx5hE3rjBClVswh
/Huv5aa++HzpKTUolXc9/8xhOY8G2gSuZ6FPjEGNo+nlqE/b14cBh3WiqzgUIkathYJbCesJbWNO
15E7vsZNhOB8PkoQalWRsEemIKnt8yjOqHdnpaWRk47VUR92KY+ItUBLxKewT8uDVSW2iiMIf/eD
VV1QkcnBdbINuK2T7f/am9W9jBcHpsus60SVG4wIm/nPjq85V/J2rwKPQXILh0x9tbXY9kJzbRCs
wPt/MGNmwVSOszcLjjgXqNzAQMa+K69ARTuOFh4SY0suEoktFt9D+NiogyR+iCwuQteF3Fru/uhe
ChFr/B+miM0kIub3GOQ8JiHDV5+x9YlZHULLUkEKFgHvu7QJPsOWMLDjLFuofsUmBBWcLAZr+RzI
d9WTWQ2FGPamNzB14K4q+urKALeIbPBHhYnkDUYZNVKhLCS8GcMg6ukdmmrLlacBcKAeI3R3cdfX
+/TAFY0dM6aNo4OkNvr1KQlKOin6A6juD+ILxaQCwcFYid1HFhU1DQo+7t3ioiKjW4wFLErt3FZy
u1EWFLCC1m7RHt7VwaVcAhkINQ4JC31qgT0JtfQa3uezNlfcsdpGdci4vpYg9WRz6OHousZ0HTDK
vtO5yg7UPSUSo7YyCLIdiwlUnJm25eoYcgdRTj6mzoKTfksH7DNxdppid+pbzuR8jq7TefdqlVcd
jxTP0f6XNeY7aPZqeQSoepH/UlkvOIzVDV7k2UAXH3NAfTdZ5j6dbCZQrhGZED0rR52I8Z70crMC
YGXz5B1GI313powvq2TLVqT56BmljjHXyj7pwIUxo+/ItpvI7hjlTsC5e3x0/4IlEw4EWazKU6KA
pId1wAFSQORcXK5A/Kic4Iltad5B9g32oMfp4IJcJOgOYetosnHv/9HX45YqA8pNp5L5IobcmvAd
WQajGq5A3W6BIpkxg8MtPQKage2aPaxqacnfTZRWEwnvOgPY/q62fEh+fzrom1SaHeTP9/TlNxxY
rGyovYBsRFuRv3croQf3SYvO8b0Q2Il4T9jcROLdxZCfXGwfd0SPOhFXBgAE7vrxv5UzbplZqPQ7
4wIiZdgS52YPZh2NBV2qWjVYsm5CrHn1oKTWBR1DZnc4i4AjwxoBPPubyd2GiC9ioYgFAo1fmhgU
8uEvGBP2omEQTKt4mKmZezCnfFs95nfQycH8iHwDy9wTtpg8jQkAv9f17RHWrPTaZgIbQ+KTbMn/
dxcB/Ng7ijO9YRlJw/vU3LSw6fS0uQoEywSadD0Zfzqd3IpnTawOEFTyyuQTuk3Fxa0qOf/FBkVq
8IG5MgtkmbCBIHD4K23lNwdFLOJjFiTFhAk1Qfaztzj6YT/zZzjWlC8hlXzJI4SOcR/bx9lHBsrk
uirnDgOGtct9mAhs5tTjPjaeJT+qNDETDWNkAzUNEEkiqxbuN6Kg4mw1qOCTrF+QZBGjlbGUEybr
ZsxCmGor3MXCx2q34qe3kIlluIDi6quejAimTok9TwMyaVVd3IRG/FN0uxPLqFHIlMNx+IG9T9Dm
RhC/hLqFbc0G46lBV9cKWvptaNDLoi9X+qnD+oa/duy+m3jO0PqVSc0GuomGCzhH4i9JneJbt4k/
E73l7EGOeBFQbUbBIMZN22eAvLfMZQNHbsGQOWfLcsEpzFwFr0Fdr6pBVWzj+N6Xe88R09m4tB5d
iTH/sabi6PmX5ZZlzeWL095WJTqvDFbEo6Yqta7f6IOd+9DLyDr9g7s0SwaLQO484bmU2bhyQ30c
XISEMilWeiJ0Xt+74IlzLgsWzSNrTpQpfPOI8ZPUdYtaE/T5ZUbxX0lU1m7CkQ8sD4Ig7o4RadiM
gqWxHvjjRM7oP9SzsD7cHuCn+RTlXwOn2nfzZHUz5hjtSPev6Pv6rjSmSRvRX9YunBuozwH4rObD
H0GVinHS/gXBKziK2DHSrEqWIf0i5FqVdx98fe4NGqVRwQVwY4v1O09RvMI2LayEsi7zM27uThSv
Wvwkk79hZNVQ3gevhc8tGdkr67Y5L7axr9DIzGKZArx23E9vSzMtDJwgCB6kcR2EZpbRGA5JIspi
rJgO7GZaHy1tYT8ZchpH6WnllDj7F2h7PEiXM3OkuKYMBAlOASMThLYH4tDQZgVhMJZrQ+AfpICC
gTUCZGJ6e/WvqTtzAL3i2C4kGg2Rj0NrOrmULsqxGTNDpyLrhW+LW52f1E3XnKrEcIHeS210ffGW
Eg58Kd2HIs7CIHYaBm7f629gwLcPveNX+2K7b65rOzEXSKlqLB2Xf2ZJ9iFQYXKLp9xn6RofOH4d
EvhqgxAG/P5hRVYpAchd1malwDzhszYv+OIJmuvhN8N45VdADd6wAusACx9Ybedrp8VvrxEhkmp1
xgSNfiZSLLWFj02hhgVvUZchtM3ylPSS74YTAPuD51s4L9nH68OXtonx2JsfoVfmDeH2QsMV5G5t
CxnIrLdqcD0YOJ9QT/5/UJrQ8hVoEuInuvJBdtOavV2rihZ1P+ooDod5Ezg+Zh78dkEetMbWDHwp
QGLKNqEzh7CzRw/IZ5rqbdXe1o0oJOsBvU1ejS4UBv+wjvAH2EmyhAZIsdOE62k20uGLyMPp+LRW
ECO43qy/7ZAzDVQZoTOYiYb+ChmNCTtT95VxdUWYKkPfYe8xXiKJphNuzlXnbcqYIiIZwvkSyI2T
6ycElP54vZqBPBMPMXWjTWxKyhT/kmfg/P7VpUEvaMLRvhORxtibI+aRY68vh7DUAp+4p+fwQeT1
93WSBjFy9Ji9k/8TNd5HLmioXbqz0gTTACRnK3ofuUS+pyowTFeFfk5Wxh4pTtsyVU1b3V7xKEdu
0AdUnyLaCCbYqvHJMQJCvyMyyhJFN6ytioEHTGBn1Vv9e0KcIICuHXaQdvR+JdFzzj2kiuBm/WOz
2zghxtEmz2qWQosvNY/SHDJ6dVhZg/cCEoW43pFIDBw7tqKZK+XqscX9jUGPJRAVTPgnQoODAMR5
mePO0m8Ij7Gt26moF5HSP3w/6SfywL5zEwGcJJEeJVKGHBH0nFdBJcWXvjp0LJVEkDjjV5QhPluM
9+VPZnCiKpxlpW/FAQpiDtjWqZRDsUqY6KRmnhbWgJ/pbCIs7fc4KjqSdLCZVlHjk7YIyEQCrcx1
gWvzaQkBfXRegsThJ7JfBhhz0nwSxpN2a0ZAut6h4MlEFDHDHs3Az/TgFwFEl/PIjOzpF201MILf
m9pAo83tJGESJVut+lZWW4gQFfVezm3fDUIeCJQO/JIx4HJKhM4nK2ENJgZYQYlvKIoYZp16cbk6
SOLUiiwz8F66ZpLGCC9VxiswsEW+NrR9UoBtiEVvlRAQjw0U/lBn/lVVXbVode1gkj8vBfcDdeG9
T3I0zTluV+V6Qqk7LqjnLmLVvQRe4U2UdajOjg9EBiJ/uR4uKPhnBiE+WdPSA7AnuKFaegpXKG3M
x2RMjjap6P3SJ21FiByMpi1G20vLgQ0EHmqO0oaEaaNnrOBvlcOJdSQL9aP8QbHjcT/0ky+BBq2Z
LNH6d6f4c+NncpLHs+07TNZTEuotaUjLKBdsdvY2wehxf3ScXx9tpMReGE/z29oO7KwE/gZ+Gnzx
GE05FalkPYzFG7QFhNovX0L1D0Mwi8vE4t4sQO25u9dlrc3SjL848Yu0ZWvzwtgAZ8oxhP/0Z8uw
nSUJfcrhWRJsxFN2jvPHF60qeDxCqinj/HFPuG5qTcc2QNQNYa0k8PNd2dYobuy07Tbk9BZ0iROI
FLQDS34JdAxv4jjwlCSUAC7NoVzBg0lnWSrpZmfEBJmoXoROXhtqWi4sjHjMVERd62AGwlpymP06
PH+47x6AxCZw5pFXp0Z5bhZe+JjoklRIoda25BH47r5vDp1E2cKlI/BU4fK73VD3QWXUscX4hPyr
w15t1w3UaOsyVtVjRubCNFwf0deof2YwKQt6rxPK1wkCoVM+zrMD/rcJqlUJtdfzuNlHg9LPvVQ5
45XEUx7RGv+F+1Ks7zkqA+d5A6QtvWAZOEcAj8Egdrnb9B4Kd9SKo7sSnvQuqdgP8D3DboQVLTbb
MFEWbg1C2XssGiJc9gv+ehDlxYCF/iyjpx6e/a0MSbs/DRcPNa55Y+t0I88sUO9GsFBeTbmVTd65
FfolQv7Nu4Q6xls4861lFAPCQcqAXfkMR3Gb3G7RBjyb4P0XGTy4ayKlBEjA4ih8c+hLuq6ZuWjA
uIY+mr4WlY3q5BlKmvkeGLab8zyURyHI6tR9FsaYYDqSllV7ldibfoo2Dayq1hrpMSYCyxmWQLrP
SkgqQbRC/vZCyT+YO+Tg32JhVUa/LQnl3NJIHYw7XQ8LHlZ2FCUOUQgVlX4mcBlcCcnztZv+CV8p
X641hfo88WEXPJCHVOAzVhOdHXjaw2z7CeAP1CKJX6SQQoErEMDtYBWsKqLr5jVDp+KV22vkJHK/
ORd1w57nynwXQcU4vU7ExA5m7cufXaEdq6CWf4A2fR9VFdQJo70pInCD2BWOD5m76QMAg2sW0b5h
VBasD3/mtRuDaAkWKi5zQvWW/NfmziGaqybV745z3ZGFW0tJg7jBo5+wfDNHsvJsZZYOzSv/hky6
d0pwM9BEhX4L42oq0jdbSJElck+RsLJQ5r0TRym5fsaR727N8sfuBEJ2uys9KSeKmFzfoPDjhQo2
9wl52dOs03izcBDqRbnvM0Rj64i/JhxcacOpqKw6xRPZx8+aJPrgkTWi0l56h5biHm9DMhLu2sNa
xrjfck6l4sJob0nZJnUWbSv0OESD6bQPh64Nnj871nHf9R+Rca7mEooXnlVZD62cywDQZ5OlhueT
14p4HswS9SP0WGkNp3XHTa1k+KLZ4SQs3IBs8uB/Bx8fyMUT5vo5eC/9ju+ZUw2XVjBC3iZcovM3
s+ISimUhEerkJ9XQbDR+y7A9sgJnVdUkvqdOQdup/B/E0ipqofwmYq4u07AjeIKxXGKxbOZvab1T
Eovly5+fKvklLIIo2aCc2MILiTsPIEY+GLr2lsCWyO4viYrWgMtFaFjQHMr0UuYiVw0nCOeXOI8l
op/Ulxn3AEeRp9zr7hs33fT27WZ7wcbc3NDcMQqDOmYtdOCi6Dyq6239NEVaP7m/pcM81IyVATFj
vd0xB+lxOEvgDSCqIg79YAGMFgUArn0w6P1G4myWR9+roYVroofRu1zKW51dEJbynv055qHaWVar
zClvlhDw2plzO889DcEQ61poMwXn+3ffFoEPV+ShFE6aDzOyz3+R/7xFaXOuuBE5tWcIFe/OD9/e
w6D/pgMtWegVSCki/5qEZfSB6zWfCrg5DuPkmZhe1oCK62ReioVKqynVHnTw1cW+o7sPFnzndjrH
uRIWk+QFAA/aUoStWb2J9698FkK6kkh5LyI2kLY7Lm6z5CJu4YyPFWsxsiO5KTe98yt1dC22Z/KP
9fKrw6aKBPw1GasF0jsxyxkWtd+c1ih02rX7lGxoOQ0XRMl6u2moAdWbTU46V75COgrC+F0qhP6x
ZFX6YTNFRbYxgUjopK5K2ufHOzOOKTfcVhV70rS7+sPFSSXzNPbYFAI/MAKS7r7oGBqS6ewAwuzk
N+4on0oapf7teIwuxXAK+p5tTNCWjjILXf4nI80cEJy/mOR3r/JOUhYOU7jRTNfsZYEFNZ3Mr+qL
XW03fU+Hc10fcj3yxpa5Wa1EDjcDJsScP9IcWwzwE5Vxkoqs38nhqZPD+NM2cggL33Zhmgaabx0a
b2pbGB76VZDYgkL55UDnKosrSZDX1Ced2brIZWgaP1KfTQKby3tbSJJsleEbZJ0/0r3MdveBhJsQ
k1Tynv0T44W8axEZ4e/Bfq1YzAd2Ml0mOwI0CSSVrnQBEWI5FyZuYOsz7D6LRw3Lm/34FRuAtUx0
BkG6di3Hohyvl4bVjZHWea1lbaWnpf98bks+BlWGu909kCGDZBKdczH/mKNSawPtwYfTFuvw7JWB
YcWFiBj3G9CkIbaOlf4KBiMJ3vRDmGnlQevwZAI2LRlcVEBC8yo3yEntnigUtdaBA7cKIDqhslkb
SaLmVQFve5NQEAtwG0/khbNHGh8asW/EtReR9UJXjUSD7je9cvpt2lYdd7KE/zypXv7RX9XumK1c
tEajbdXZzgzISoU+O5KGGyDDsfrXncGuJWi/DNm/wGUJgjpHLchRRZQRc8cBCEvSLyrAzvqlbCNd
a2OmL+yX8MeFsfwSSSrr0KeW9j+WfA6eZk3QfaRmUNwjK8f7ikn00EBnwlJ6UkWDW/Enjysr7jgY
i5HRAkBCXpRXarNMKv+Dn0JOG+2wH/wLrvho8XJeITdtIQHu9y5XtClirBkTka91hCtUeLPtg6mp
Jr8Wi6P3CRi7O5eDGLA10A53IhZMej4vxi8zvxH254pfvED6Ap7zLoRb2+oEiIVyZ7VyRzF7WuQb
teAaTwLh8Gc6BMO4PrqaRNrH5x5V3pdD/yR2eyAx9vy0UzMwYlxkdX6EmBbApIBs/k834alrNYEf
kYQgj9i1Xvjlcbp5awcnD8D+JeJAHDotjt8CKv3Q4LxRrH6+Ozdw/M/p/lsPhk1BUkF5Wl18hKLX
AqSuPcVOUGIAQIhPwvmkAAsqA+mOMpVf7qecTcU9WLBuQE6SuGNNQPg03uBrTeeLWfe2EB+Taf24
XWsTOrnYYhvrRkDsaONgqXKrBpuaKN9ri73CnDcBHiDz8HRh3BFCgdwNA878zK442Yb0AsfqhLpQ
3xIOXIqp3cKrV/Tq1nN30UfNNdMDGUdYPVqn8wPQo4UdvxA1fJeOGWwsQFFqCie1U2BsjQB1PaR5
jVb2ECOqSfj1wsi8lRtr+j7AMYcGRXI6KOeE/SpfB+LVZZ1gn02YVwbIrZJLjWzSrq6aZprj8Yjt
cMo4tS31hK39DIvYuNCDLluRovUGEw7Aci58bS5BiD06dRLZJbaU9DMNrMElDTvisHzHjBtQyxgr
DrHY4pgA+RL28HFHHGgflzfgEwVwuyh8qS0SXs0BcVgaGBbqcZCYXcQfcfpuTaCG20RQHSwZC0ct
JNMyL5NPguqsi8nNGnLZHfQSUumlF80WLgLmBjYhADHZ4LWHwTLD4ZlPnpBOtZqJ1COHPKgQl0cI
t1CE6qMmom+DGjpfAv+VDIFXs7RVwItI1DrSGWAxxaEvoDqxWBdqnaMPJMhHeTivhWQuipBlZQlE
C2fz95u+iPyz+R8OzVId1wgob0fXgx0XvTjfr9eqGA9N1YrYoXkLvx55wBNExwb+Z9xUUa0zWlD9
tRF9TbGisXSs3d0iVIND8GSfpAxjfLX/7ChPVSek3fflLizGpZbOyy6jpTlxGW61mZltczdFs+lb
2KxX5WPOaFniE33Uq6t9O/7+uOKJ2XiJJtTlGzt6YrFe6n3z/FjVvb3Ysh3VrLZ2VuDD3CbUFToM
nKQp4VuaB119Pk2j+ov7GXzzFvPV+Unk+3Q+l3efIJK0Vu3rWERHwdWMkinPn+VKpLo5XvP8ASkp
+KuDBDbSrJhYB8yXH7h//+mfcXd3DlOWMSKIvu/wpnkc/D3YzE77RniJFDK5LXhGp4eEf0SEOgXq
nzMIDKPHjnkcksv8WgHQ8993dzLojPN2gRFYEQMKzIaLPxHxhTqhflV16UFWERGIsWYy7KX/gX7B
mO0ky3DYl0i52CxtyuLBcDIIbttowzHQC6njbQxg8PljKoIN/WM0uDyCDhDFX8guu67WOAD+EGql
MIPpy+rov0U+LYuA65zwwkPj2OvkasPa3l5xV5C6ghalY9ClaJNRShMuoGK4PVfcXEkLVFceUKUP
+wUfHOWYTEyilpn/RMA47ogPG69pfWPwAI563dxNifDJC8yJpcYDVyJ6PWnIbSFv0p5I4X8FyRxR
I5mmO+qgJD40QSU/ss3Ru9HQd5P/b/0q1xeMV48kIeXxKSzCwQxPAzs9ums4Jgl7fERSj08dtJiF
wIHUCsHzom2//Bu755KfiqLkp35ZvXNQEzUrClzY1JANMHC1NqjsyvEc7S8f2wakygZQa6Pgw7xE
k5nzyxtC2bR5jV7o1RG9bWU1HeGi9eXr5hki62aoKC5avvjxk31TOb79q0DXw3ZRSmWsciC8XnHp
t8oXzl6BL1BkkqjI2Z3bRpi/wFj2OHW1rsp80SILf8sme6f3wQiOe8gqq8W0LMCowlXBK+/ntPZp
hnZbEw04S/JOqLXX1iJTV+jUaFBpv7r5TM0JKemAvE1Gj0FLY1poUnWiUKuuQGTM9y7NzVMPU2q4
xjXLN6YQ36Z+KVMwGlL3HFrFBkmcJDILvmA5XI9e54z6QDMN/GYAUfz1NcI0VN0rCvde3ZVYS/mc
AJStfudJASnL3U2IBBBKbvgu9oRzt9aARc+N3Gyo4wZ3lOwg+Z243wuEtJn0Q2N2+ZeQwbTFrTy/
mJyUWanxzBGqcCSu4IhNDYWMqTXOGXMgFBgybEV+F3wq1uk6gytg33URqblfFtiGlVAHCu2cLU6K
/mUr4Hz53Z8Wujg8wQRWRcNL0AQyDEvbHJcm4VY7cxDyps0QdONalgjTQP2LYSdb+hROLdNqR1re
ZunH/aJcg8Nw0o51qJAh/O2YxcnufoJwiwnwcx+oEsfhVhaA+ux/KpWbGbiq12KrsxlNnNWLpieF
Dm0kbMJs4uNYniryquPhyrnyfK9LWGrFE1fDUyCyrLk1Of4emHM3qPI6Pex2YhRGzw75DIjyZVkI
3Bx1YmB/xcM5IBVErlMXkTgmGdGZSv6fbL7mAkusmQgRh7r3Met48qu+b4PjYskWSr9Z1K6jj/Az
OGgJ6TrwnvWdcnuv/+GsWokbj1l1QSSS2k4taxxVn6RVf5vQlbPTCgF9nFatJX6AZAf4NojnQzTU
T2fR1JiyHKXxHafbeFMzMMjfoHXkoGPgJlfcqR2wxQEutJxMOS1d+gXhyKLGxPfHA1UpmS8GUcAt
tqamUpkcApfbdmD52aBnWUdGC/awwWOiP93YwTeBFUFa17a19bK2R4zIT8814YQwNO3UTiP3k0my
utLUSe4SpwMq1Pvv4HDeYUHwFX3GqJeIWx9anjjOIhD9N0RCrHvZOygb5YPEVVD+ROA3t60dJGDA
4udIbHUkKSUhYqGNpXdFohxhxN4y5MSwFYT/GV4MwjlUKHBIrUssLqtopd5e11T4vfUHAt5dn5sk
M0LdWhC0UHS2zJDCHNXwhqPHttC99M5briXhpCY0Wqm7Ro1UF/X730k1SrzgFgu+7O8WZo92yF+3
v38jrpWOuHz/7ZpqhUrQxeqbplAm88+6QTgqmVevg97NuF6vYFjIWkV2cmHWKY2thCH3wHq4uo4T
wHYidorlo/BttWAR8EKC7vWZfWvhepfVRjkG0Ruf1CGcp45QmFUD85PA7CEGsg+fgyO0pIDKbzGk
O9Mf5nbLWdmBJTlyWXSr4ux6wNMJd6dYtbWNNkEYy3GMUTb8qxgWmv3EN2hKBRlYin0O3cpMVlNE
CWrS9YrK/oGQ6Q+yM3dqD6ki2tOUXFdv4ISMX9cuZlEIurOcPnn94OG7/JNaS8aceAt3kCM6rfig
Zq6+44/s4SBg2t+OOK2fN+6Y72J9YMqT51oNa1aJ8vb0u1XY4jQXlOC8p1hP1I+DsVrd+QmrKYoa
+o8x/dYXOiA5WXewTdSNf/VZ1zWrb6a0EjPcIRTLdM1sV/oTTJRyJ30pZyPTL2i//KDqInD8vHjs
MjU2F9UMeehnO6Ev4LpgyzSwQcZHqY1Ex7+Opb93TypDvA1Bm0+pioHjulmKPUqMZZ/Qohe+zeG/
398X8kacp5Pp/J0OXagrtHUmnQMaLAGIIcPO4BdPFkwo3DzuopWbJO9eKDscEbGFUTPPq/BCWnjX
UO6/z62C0FTk5nqIOENeuyvadN59PwvklO7hlHX5WNXcFSfkurgkS7DEc8W/BvQst79XzEdLP/Jn
p8eXfTBFO+RfbAFLQo8IQLqZ7lbMh9aN3wdl50X2Bu5PMwAq0/gx+ZyJbjxkAnDzYAEQkLsMLl34
0e9q1HVb0s2OdhUiAio0EASsg0QTeEMxTIehS/JhZ8MBxIgc7NVPvW/fqrhZVOx4DKBaSU3i/RxA
V+aDulGr29K77BkE/PIuOiCY5wuknSHPCWoFQpbkoqQhXulvujGzn0QOGekezul4b2kO8ZqS3oMh
gYo31pOxRLxJENG/4TvFyhh9uigE5SDaYgkcqqCxL8Q6FjSabQ5QQ9MSGyCBayHeOhRxNIXQtdnF
CjlXP7KfTS88V3SC8mm1uL9jBJofCV95b/SAfXRjYBcxEtLbLN4uHPLLj0T1O7jz9CbKF8s41o6J
YR5LoV0e5Z9LCWKY9azEqTLsoTCKgL6psVgMXj22LNUZjyDnwemXdOxUpFbCXDLY03KiOHyD43hk
XUSNrlFTSH3BOZUv4cPwTdwUk6/XEIxfxCm5NNl6Ql+Z3vYF5PhCE6gMhy0E8Wowf1hm9jlrU/kL
YMXUFMcMFFlQSYGWcD+28SMaqXOZwUo1jsLc7uoeO8hDjrRhGe/NUR6m1fqX5wN0jICDjVBhyM6n
xxHGfISMTQZYdBRN4SDcS9J0Q4CTxv1nunDa/rWNKqTs+0uEuR8le+4berY5Xt3nRASWLMVyqve0
ff7kiEwqbfTDgDJKJQ4YmeRBTCFd94HKCiGyqwLmcO873XMyl3j09NixcESDghiO5I6tyDR0vCpJ
OCil+3xdPkXoLVF8niyGIwEXD2i4a6yGQfTpTQJ1hS5LOQCmfhKOQ1Rfg5MpcWd424bZlqKJkOF3
6ANryUc2rs5q0BKHTyiNGaRtoyyKn5fYsMSJNAkAqkR7EiAEF2V5nryNWExEQzIPqGdMAnPSpEhV
4ZutU/P84cqi+4Ieu3dd5HtuvWv6SVhpnMQJ5O2cnRCWOV2tOFiiKYwRmPYQfq5tYMvwJ5Mim2J3
iNy8Y3iwjrhwhsX/lxoohEj2lBovKXqpKt8BQkFuXw5YMaJrZ6fp7p7yDdURB4+Crz7nptpxu5Uy
4Ji1+lWP8TkT0yuy2OnPZ5VkaPiEpOD+M3ww9Ed5z6ZpJzx3StOkpqyNYMP39Gfhh+mushvO+cVy
p5zaXnoDv3cieEMJdlY2UEncl//r94ZvmMpsSVmuOqW4x1gYFvjMW+Pz/FSy78xEwzj9zgEVpj4a
WTObQZZymdm9od4mnvhfrk44B5i33JUfnHMcAQfFm4WYUZGEu2/mIQjpLk2iG+uREb5UzeoyXGJN
FbEhh14Lab87VDKnIFShIGx9m7CMMuD1rWTb5l1sVNFRZLxgmKc+UU8lvcLLPDYGPTjahW38aThB
2mitWbklQsI/NUXTtRldAc6VrrMWoQQOe2wj9ltl7hzYAWfYc9L086xa02fQXzoDwUHZClQUbD5G
J9LhOJ84IN2Mr+kxaYiOd1ntRSpt9AVX8xgo3P5T/XpmgbdOZqYIxfSJt+PuiChLIN6t2YEvCNHB
mmkdQoSxnQEzvAyCl76U/Lg9TwQU9AF8R4xWuW1csSoiai9qc0t1WpYY7fMfKv4t7pUrXHew9pZq
2csjrsyyheeglw10y3TUBcJVZfnmbNrlON4NX6L4vbXY47E3jyRk+f4WA1ZW7Lf1BueuhyQE0CGp
6kpcterKheYqDEEkTSRrUx9XMtpg2w6KxXBJGD1xO0DUUlhEjC6UTvQcS9bsm4iJvHmpKSrx54ZC
hJoPUf12tQXJYOvP60dD1ZaUi1/XvBBVaQLZ/BsY0JzluBTzhz2RgYZp8dWfDjugXhYCU/VxVX26
xzNMH028Bs8bZ9x/+IsZUv1NoU1LrBKm6q2ZRRozmDv6gY/a6oG3CIh0LuWS/OzslixrF5fW08qL
jlWLxSHGvFAx/bXZYRCEjBRlEJGoa/N0PnlAhNe2HVYw9tPP2mabGcv7otg7Teo60jeXvfubcIrA
OvtmNnREHlAtOh1CD2yM3/L4aPGwU1gunQjgY3Fa0JLC2PvIxVqd2djSqPB/rY5V/285UBNulOrr
7vRSs1iSAPmdAOxr2cFOEnrN9vZ9LBvugJVdu73yBTCjzj07VUINzEAto+TDGjRh/rXzgr0MNrIW
ls+hdjml2L3QeAucdAlncHUsupJwXJUi5MED/A+yxcPoDZifs9QG/iMCy+mbjuDgrhT6B0hINa46
tNAg+UsnoND1Vp0qgbH2kAIGisCBfnpBwJyjyRfvS9AzCNptZ90i9XsC8+05hEUu9/sHS7J941U7
3haxzWk3TAI4kUM/+3Zhf/4p0ffRuIQMSiCw38t3/KJns36oIJ30lq+LGjI+aiv8qDGiuTrMFB6p
26MXTDGy//MpXCeQns3MdyZn16iL+pxlEHpDI9Dvg1WKgqC3KE/wxR+RHrJpREuHXxvWttHvDaS+
q+UoDvIzpV6b/9dn8udjCDQ9PZgRlRJ4oel1IeqrU8pIUJOXLtM6dyXJArmqOgpFqhHry+CIrJ4w
bUZ6+unngWPRQAaworKDC6kKqqq2WAfdhePFT0OnDvqROWUfWJZSFY0lmRLXF9POg3oMnw08Vi6B
ordvLwUukpIlCf9yOB1rCNn9ugllpDqoxbFVWSbXCO5M06ZWuFjnMWtFIvKxIc5NTQFO+Cy4wJMr
jTQ/F/wb+XjkujHBvRlZC/4+KecfVmE64gxDDtYQ3yM1arx29pvnr4LMyFbU8mQHz6PKW8bjJgMc
EQY0Lzzt4e9PX6H/XslRDfJyH9yfzIaA7Qjq1LWgSLtKb6GqSmCxWdEa3NkIqimlnlKsAZT8QKkF
vPVbWeFikoQicHtY8f1fJoB2xasoUEbrhe1PNQdO4P3AMNALlWCxk4/tC2/AmD2vyMfigyZPOmzm
A8bBGOptTAmkRLTyQ0B3Zm9tDGYiHQL+2bL4iwAbcIMrARf5IoB3FrukMQ3O40nNDOPrB89rbEwz
x3w8pAQo13TUSzc0jfgb/Gj+yriexV0gHqdRKoyrgBI7RG8zIFLVMLzoEIxslA7/LIIIzSLFa9Pp
OLblEoLcUnG6aPLqUmBmDfIw6+JfvrHk1Il4/dIlONsYFalcwV5btpm8pSWtDssnHigWUGxXvAG5
h43Xx09h+XpCj2Sic3dL1VvB2i5PoUUm62qplBLRauKgr/3R+7WhtlqjdbrRZ7LsBZxsXbiWtRzI
DZ6eNOREGyHfL0Ny/VAFJXj5yiJ9/CbzkI0eFA/OjxdJ6vzY/yZpuFIyxt0+l8i6PY0sTmgw7YMm
NmuSJwSWXIPhPjjtD6uHfQDM0Ofa56fvJ2Us7MJVWGYP51wj4SOIwolMz9WaOTo2t+C30zUSU0/m
Chh4fYWgElbSJDADdeE+xSVu9/mxrkXlywHM0QjUqe8b6vGIOttGKW8LtZxh3qHHDwoALnwq99as
NTDiM9XJfGWWk4Cq6SRs/itctZCnRm2nf8zvM1GrLnnL4oYRgx1lvCdNPLf9ckpf1R/2iZOBcdM0
FrYcYLptwmxdWs4ukZh9sMPmV9HL1gMASBPT3eRsM7mu40ySbcTJVOoHwbM4INShvJdeg1g0Cc+8
dX796lWldVkoRHz9uG0yRHZ2eA11mTCDquurj/6tc9V4qyZ8LCls8mrsZwyNBEkEXpMfXx9TIXUS
XoD240RwDTp+JCLwqerMfJS/ZZardvKxoGIA2nBenl7UK6Rjczf4EPQ/f5SH4KqF/axPJz+chlmh
zaEQ8MlDCgz5hxjf+bbTlloPON4kZlq+KAIFWr0SDPVwE3NRR51R93PoousZ7Y9UUuF9WbMFLgEi
9fGeQJOWanhIYLMLT3qD/24Q8VBrEVMFV7VDJ65HQZi0t+JuSN1v6c3BbsWVzcqUqdEXD+PAPSgB
4v8HUXHeGk+O3hnNGxRQnlEKJnFYg3QK/yyDE4kujcAUI0Yd13JYRglmOWzzAy9zqJNQ81j7kaw+
bDpbZac76JEB+PCK0Xn8t/lV/xpt81FZZ7ofcjTqxqgWUpoqJDp8qYDx4/2TRv+YJBE/DjkuO4pS
qnMowXMXxtctp6LhPKINJxL8aq0Ex1D4NeCQAAs1mCZKlEtu8q28P8EhoccrIsuW1pxIPNC3UkVj
SJF13GNYa/CtMvDEDdi6LPNO+gDJ9zz8B+QjwgRWiiKjuEes4bXPZGsMCJs4XgieNQ+Vc+XZzgtD
cG+HYC1KA5nwurfKSJRVhjKgLvFMbhOab86XefYYBy0ji1ieazrA+uROU26VkGeh68BcL3bjnv6F
GlyQ/V6s3dpHUZkiGukgCWeMKFpNtVRNiSE3O7YjhKsXI1S9AZXcGsdU0YJitMPUJttgCSRnliqd
ZTRKpEUef/8YVnbBJSuNrDSkGqnfCFxn6102OQnyHGSQ1eIPpK/oOO6Bkn9oHz2b4sKJom4P8fSd
iaoubCB+K+UKCW9OJ8fMRP0c2EsASUKfQyuOBWkpXENrLymjJNC+apNv8H6TlgS2i37Dl549sQNz
Jxnw45jRmo9UgmnVZka08ZpMWHmbJbKZFeKVyTZH6gxa0vtPX7tWrrTGI5fvUSrEPAmQC0vGLhQn
wYRpd0gtYUeWU3YCBKGhpnBu5Nq6WsSdILNvvuL3bTUCiZWcui0U/XMr+01WirK1g9hy/raN10fT
W6S2LMIrq1DWWAYwFKpcw6iRKy/kbmwJB8Oo0vgsbCQjJk7ImXGIOrjQYoTLzpvjzkTfNYOJohvh
wWSAlaPJZ46pZK6k+96I0sAxbgFN+erj5c96n3SjW6JtHe4qks5bmiQvOvzAEoY+1diFO1s/IVnK
R/jF933m/DtCmlBwLzOqLMvO2EvOTwL1k0FUbgqPU17iCxh9QLGMmOh2N3IKLMiKDNd8YvTr8F5c
RN567VtjcAv3c3jTs1gZWosy4dqXX8rsI1sbrU0MUmo+Sj/vzV60rWPWqs4xVJDc8Hbpn1Itw5XE
FlSQ3y7fL5XdcbmpH2u2rjGy9d8bjKYa1BRntqRdg2zUemG/sswgqbtJyu1Eu5lFnIj/LhS0ApQ2
hEKto+N0RrH37z/2JW2/Q1wJjB3yVVV5OdeoxcgQ3snlKu1+96zOjVeME2yn00DJsaB6eGgMRF77
gv7T8HW7k+uev1vMutKSB2oFrzQ/J59J4Q80cEl8ncYbCK+oUB3ux5znR0diQfq4/OiB9Zi0xR96
3Nu+EOCyt/5QJvZirkB9tWQlcoQSvxy93GExnwKoPwG2NsXN4vaBo9fSCi12KlUiHE8NEK0NWmg4
dvYay7lZJZwmq67mdRLHmVQ7TVvSHorB67F3wxVnS0Tu/S4keDAafwfteT3LLOB82N5qQbT2aLMy
Y5A8RfLUYtf89+JuM6xtkonnfWzsJzS8O74zRNnXDLoOxOb5vtc7dfVjPv8xWf2M77xUHm0moHh8
3cm10d2DDeSzDjM7oT6mfhw5XpEtFvUZh01wNcnJk6IHoPOjcVxP8DgemhF7viRSeexwa50nY/95
8eqB0cmMFLgh2Y2jP/yCLIZ5C3YIMWaiSPRV9Ft1AZncsHRXhRVKZIFQR1vH6yUpRT3NA7vr0QZ8
w73KkuR0xMuEdpyPvoZ7r9PuqXvCtO8oHvmmTVLnj4ppfS59+5hRYibQzw1SNqoArBIQ3cafPHzA
O/VFgTIcwZTXHlSPK0eTphBe4SzwibhHiJ34IFCSNuclaw1+Qb7618ONgyNAK2z6bkMHrYWrrcsY
w+NY53HU3UJQKsJiJWnqouJRvcJCvrRjXkzHzInB4gUy+Zbx5Sjk/xI4m4HI5H5OuDQgfTcB7QfV
cZrIWD8Yor1mX/oI0DXhscVjS1GARjRi7oF+bCPLqvzU+/2X5rgaUBorynjHDjJtOlb7AcxbecIT
9nka38t3MZKzpFybwFh/A3xJhbF5f75L/3SAYAbxwQg9NysK7B4C+idqXMlGXLVakkgZRlbFcXRW
HaJvhStV0LMWzw4HJ2s343jPoovvpbYiij0IhQBgHYFR+6dDQYhSZ5ADhuS79vCIrbm/BzzfB2CH
5QR75NG12xbJn7t7/bKcvqrnUVq7jP4WmLztXgJJhxD6AQ4vYzMx33IFwFu7fUWaErzVRfxhhO2r
lJcLikJVEqmwnH8fhaEt4TFZxJFX9nObcq4tTUaZ01rmNnlt+nxomSu+EFbHkiqKqtQ/+Zr5EyGv
kvuuKcSW492lzxVFba3sXQ1akCbLIjeZqot1vfs1XBkHpx83Eq9riu5piY/6hJbntBjwNc4tu4dp
5rX9WHmVN3SCnHVyRo3Lweczq/pk4Gv/3YqP50Au0h6LFEdY/7Xw1nX5jumIuBV+FQs99UHpeIg+
6I1rkCiFEREKYl7PUaO7Jpz2u7Zld9Qgp7c9JhJEi6HqIZpOE485U3uYtJAIi4eOAwmQ3Pe7bdsH
PrVEsBPaqlP4OZO5PfLXoKoLvE3+FWCEd2PgUy+wtw30l2HUgMyQPUQgk43ZFAqBCWyBwKQr+KqX
gw/jjSL7yu2+lkfHK+ZcKuS5cj6kRbY9GjznutfTlChBoDuqxeaHqxbOmr+eN+WdtXDYAqxlpYEL
g+vqyv1dKuoFiorJaJkVs5TWDDMbkelCIBBttlBgFfcV76zKgt0mstrrk46lOA49wliko/Suggey
VcdpEi+R6EmjPWaOiWpt/21PSlpuFQdtjKoKbK1l49hiBfR3HB+SbmF3Xdcy0TxL7xzFWnppJyBf
AMpELEUX5FHqoBoTFp0wUxjYAbxeyXWT3VMS1cIo9DsR2/PWtUXaZh6AJIwRNPN6i4Fy4g02I6+o
C/TGnOeTQuhXlO9PmHT1RKoT5TaVbJzK2qLkZTcACJToai8psNk9opSxHZ+wP2DYA9YmIlPH+6gC
Mus1B6iGdf902/WT5j/9KBXUEmka4a/cIKBjTbdN1jwEWXa5zj/EU6YTLTY51Hx8Igx9RoyZAKaJ
bJPPf0PCAeZ4aWsP4UiLWBGGeWSQ4xqtz5Gsp/SpVg8SFroiKWvkPTi2j3DR29J2NRgIaVqKMFf+
WH6NLYcCqvSuCs5efB9Sj39eXlGXEjzZj9eH/0LK7C2zPxnmB5jrrFHbCuV8z/SJAwIS2DmFCNwO
6Yr2tswqYNk/IOWEfmeryujsNY+Ykvsjvc7N1AwG+28r5RSRxcQesS8I294I+wMvTH/dpg4cODv2
zxSDH7f27oA99L0ZaeeBy+Y5N41z/ciGCrN01tUGNvXDLIY6Vm19VLKUBwiqoAG1HN+ZnTG6nuVS
tQlarqWJjjCMyhmtz8XWcdkUS7qiyap9JYBUvsBfF36s8J5tNopAT5T0kBTb7N+4wzp8BE730lC1
Ah1JBJguFsD0rUePsoMmMCm3K03XD3y3VZExvXQcQmlV4zZSLHBButqchS1XI0ZbmpwxNw5zGzMp
G64nmrfBPI/55/e/lS89wbtgGcZy7lRibvpUFGeqCyRVpzpetMkiyycDYa1xMxCLUgSodY3KynyY
hsqy2p4c8p67fDBvHm6fNpfNJDIYlEekLbjStDmOhu5wgGdMTBU81sjSA1KgDPIFEMj6XmBahTfg
LYAMUnTGmjK+4q1Immj4v6DpWvggkXf9xdFMXvrcpgFHAmc3EZS4hJfqGk9Rkco949tFYhNvJrKQ
cXYOTdL9DTnxnKQSxIN+lMBGer+AcqaRhqkOtRxxDTyta6Bfrjg9EMTEfOiAwXs9I99iBKa/LJXM
LLU4cDNg1mfm2CxRVSVxjMF5uaByd/N35dKBHvTi5gz/xi9ikVuYirYVoVA19vtjvKcgyiy/eycK
kfntY/1WLtU+rVILUc6WmU9fui/Jy58icngDoElqOlCY8zfbJCh7mAvoWUlNeHbVhM8N+cnTdzsA
sXn6DqnI2RgtNmMK54vCZJiaPCVkupOAM0eYZeYDJKGbfB6ADMwjTh8E9k8XL10qWxlJF+amGcwa
NSX5thyaG5B8FOugegVX9gNSlR27ou4RvNbKZSorQ2ev15rPkt3yh6Bs1zi4Leov+SuYVUQW2Tqd
0AFUzHnyJj4AEZPDpKGCRnUsXNXvgWXBUf+YWleuIO9Y88za9w+uwPgHt3iB5HSSEcLG0nUcB+eM
Ki5xRUUy/XlNiK3eVcj2sAuQeq3Y+GlYF/UdbDih1EovInTb6EDTnBBtxDkMlqsj1XNbl/uZg8ET
eRvBw5McSxlmovl9Fp55V6js/YrQml4XuZYof57FeEZM3J0xkhVNphZDiu8F7BHpmn/CtK/B3eJ5
av1XB94f6PCSxLQZnDaD2lcazzucOeoWwax+3WPBjJG9AfbY6dCYgurg7ovxwUj1uCbH9VIrjbKh
2hXsD1OrfJsDvhQ4bKmRJzl87O5v9CBKuBPnKKHk8sqq8sU4ai+vNUGaUhfJTwIy4AQGBvqd6MY1
6tHDej5jlyRYUS3PRHdSPsmeUPPVxP0VyMqy42Wkt6ZJubkHfv/Vmzi1lihL9SidStgnKVNKVrlF
dJIe6aWCnNVE474XQk4zX5n0H9xFigR8rw/fbLk+PAv2pdOo7+POENwvkt2gWN5wb9Gvu5UWzH0D
q97QwfVvh4gz3fskEiimGbbO2mPdCgoG3gKAGdK3pdV4fv8MGAnU2CSOyNYdnVIdWdrDSzItQjVs
mybmz6Dpppo4ieAvKKH1QSTzt6DTpMKi6h+lrsenvG8+XVIV/h/Rk6zOSzebl5M/1u2Tw/vr3jW8
puzDD7p75BYw5oI1y5AruLg7GRhNMxhKhYALBkwrDGAuwQNde9igT31p20ziiwoejttDl33NEqcf
CVO4OWIr0PFOsA6uhePHgbHtTsT0PKO0VQsw8t6r7ASonhxgwrigqeiBBqz+YZIley3uryp3EqBW
gOdpAAOyMJ7PaPwYiXqnaS4/dn6QBmlbeSlC/ZL1c8pqFpzTcLUu1yq4Q1s+HfeCG7w9xG6+GQXq
p3fME+uh7RdxQRJ8kIfcBEsCwgr7dE5byEpOw513WcIvAx9ImBsVUJkae6MFTHrk5cszCLN1zqY6
ihuFY1Msmg8R90mZDEEjYxs+x6OcQ+xKV3fFEVpH2vPOS5y4LvpcrqL6bPQhIejJIBlmWKk/5rxV
KpVXWGwvcVjYa8kJr+WA0b3uQQwXw9iMIj+mCKGNq+Sh0jreWZJGAupRCtCqFSnCby46o6Gjdubu
QlG90MKVsUFSwovY9/0ielAWZEHDubZnDqM6ku7w+CWkh+KN8PI43ND7ZH4QmjuPVC7rwznTyODm
dtldun8OkTlb2mclXfZMBAScP3bn8jZbxAP7FAHrTQhXSK/j248cC9OFOKIrB6qF/eBvoCVUSqV2
nckWKUFyoeBi6xgaqKS8rqEVPKjiT5F6EgOCgUC74J3lV2iyP4os6XnKIM4RJup5VHbamPRM1p5G
T2SrKOXp4BLsi+YccCB1Ag6FcG+6qjROo+h5wxsiqJ5N2QS07jThzrRry6eBnenE25UYWyJ0sCZS
V1BHERmTnOR1wYDVUbcMJQrPz/0fgDrjmDEgYgodaIFvIvB86IXnAdV99/vzJw1qn5iJ6sDI6OxG
ex3ZsRXW+5kuIfapzqA3PtfH5NdJIZTUuCoWcJyUbyoL8EyVI6xMm++Jx56VY0GDQXwYmVIS/xtI
8AWaGwmexhcYHkVzE/YmYQ6nUvo8Ha2+6VNZh+lzVE4Bhh0ytFX8sxx33TuTpqqcHk9wOGrbNC8c
FjPCoLgIlu/cfwLkaY/hQB1HsCMQqZ5aKaETHriIiryzgjqeSY4tytvAvgZYMU4iL0qOq0S1Oq4h
olW3wcrFFzICD5rgZJXaPTFANlH/CxTbdqOPR3vKyKXyISa5OWwsz74qVr4pBOQc6sHKMOMBCpLs
kwbbIUdxl+Bcj+vOTXK7HuUm2/5ZaHjm+b/kda4zX1vn6YHjyB5mnAw5VkcQrMDeg3YDt0jlFmky
oMj4BsPE2+26b2wSVNCHKLz8QFvuO8XOEEHR9ISdarDxXLVyqz9QhyyyS8ExhXlymGa9hmsr0s0i
MeevKJxzZh51J8+uqfwm0v+r5OUYAWPmeLFtQK88RFvBgITIgY93/nlcLshfElfIM6DhI+Dte1df
RIA4Wmx6uUV03fFQaXgpv9hcbhsXNJPcviuKEK5kCw4ulLbwBQoB3aZW0EJEdXUnC5PyxGGQh5eT
0y2FR6BCFCMV9B3BVaKA2jfGfbFKzpAUP/0J7JxWsRdx3F09UK4cyW0gGsdJvZ9ChV2+aeJ6BwF8
+hMFNAEg0bZy3XdNP8K9jrr5TO7rsvhHVhkEXMpAhpmsoDsCo+tdAYzfGyw4vRZ1JA83xLZ+EgB5
Wkcg++7wMXGlg7xO87Be/owkF1Sqk4LHCh2tC3dzjzf0pIFe1AiQ4dxDx8TJz9WYA5Nd9uwUxLGe
s2LcU+UwaFX0Y4rIEJpp59oGw5iWUcEd6kQwRwKz+CzOdKxK7+fDdPuP+lXixnE324mI+EcZNINz
XOTe6+x1jn6sfuhZAtRokRDf5CZ+ZfJv2/oQ37Q3swVP2DIzliAPtp7Emh+Cd/SehVUu/AKmW1M8
l4w1yO0qtqRESMI5DPo0GXpaoeZBZIMDAC4ZSJ3fsQWhoiXWoDrzpuAd4/j+ql8fpGbnhQ/PMDR8
CDVIpFmyxjwHKye5SMD9cMPP3mA1ec9KcxM6cR3Ulsk47kkfK7ZZif5yZGtwrEiNLis3uHZgPXW6
SsLYDDHF9hmJjEuiWAvb1YyqiaI9Vu3sKFUiYg9X3DXYQiyWoNax3eKq55xmufXry1H9jxvHLNlS
P321vejQLg6hLd4PKUQvzlHW/hBALGpOBSkN2H/zI7p0xQzf+Xxr2aiI5/lfdU3A3r/vqATlxsxK
I0zk9vz15YcNvYFAH1XuVdH3ZLlrKhuan3rkDA80Q4SBN4t3L/jv2NXRhQkyJkmSZOq2x3n/uGp1
7aV6FRfm53Ynuk6vy/dTGGPiQdU/rCXpmOl5FEL/xYFAjtlmAn8v9mvWsnysqkmVBnGWRepYOcCs
PuG4cAE5f00JIv3gFacfWEVJCu+JDJl0wlAf6a7NrnjiuMmT6/J6K25YnVRkN9fKdMQ12hP7KfEb
waoEMeoM1AGvKdeqsgsYLJ7uEbmBxaC0vNdHRdrYgP2S2z0Q1Fo7Tz+BU7YH079WIw4lwqQsVDvx
mIAdRdqqIgqbnZSWmmSGPCJQNmLKMIQZ6Sw3wNapyqw6fzN1j1tm3vKNoLXtr4H0QBM1ydu+1LTW
hZybGfgFvf1MaNDx1ZLKC6kw7t7baabqu0FT4IZDZ68laryHp0lJ9nEhKD8awBQgyvqZnvj/JN56
YER3lfmipmnGxk/sYUVqye+VwtiLX7WxFAPu7W9vNnTTK+xlJvnkqYHQuf7CsE7EazvdxKl3DlfH
333IUktwTbcW8cb/wWTZafhNhrwV3q97Jbmrpe5b3Im56uqB/N+bil028zh9GXM9fkUZA3ooDNET
VM8pimRAf0X3BeXb5wnYDoUdYLG0JbJdY5wKPUAFwyxKvIUBlEGimh8BJ0FfywiNUr5iXeLvjET6
IIza0r7xgRXYBrr4OmY1Q9YvGcTNEevfL0ZmMqLafZWNOpbSvNvCb/Z2SPKWdSGDO9JiwKW7gqv7
2VsMYXvisaBhftQc+pXc8csBXeJO0W5aGHRwBWozyYgD3uH4JasRfJE2Ur4ExlwdYBsQSfW+onk5
gttx1z7s3IQioMccXodw80p/8TDj67I4j5mWtZptJsCX2F2Mjxl47oCjAX/Hd3YKluQ3hOnmV3o2
uAzznxAdCq5i/VTMUEjcq/Fx6PhxftnwDQRnmQLrnjqqlBKhTu5DFzXOUgDCtBtkZm4A76XXtn4d
kvI3H+qQTBWXJ9pA1oIc0hXJLsvZyTBpeBXuANtrUOgeZ45d2EpzkyR6vNC6ZNpCiA0EM9riHLoV
UsOZ/Gl+GIjPdYRyf/gG7xjxzwR4rX0PyIhBc/FLN3REnNOvtUvVmbmn/0qTYOuRJxSqAIge8DqV
PzP9B8BRhcmS15X04YyO/B626lJH1PtlJ9mqO2rKfwSf1b9JIR/Ll0U23ABct/bBTY0mJKWaInVH
jgSfhvHE+rY2IZR/rS1+FOIDxeQBtnLcaHnyFq06w20CL7X9zHnOD9ZecomzwTC+tNnni0DilKs8
+Q87sXxoypgKV1TXPOTG6IsdFQmunSMPADlPNOjwY+gDtu76pxjZ193vDinQ5fV/w8HmkQuPyl+q
fRZwy6CQuiI9VjL1AeP9NWTIp58RjxOwdFQg8OznjEfCOxJe5nYIDitqgu59+TmPG3NqLvbruBOI
WgD9vTiqOhVWBAG/zOPNHoxhKtVqOnI9waxE5F3Igzj5aFIA3Lre2is2Lt/Uat/53y8qvvtlJeEV
htKNX8Bot1ZCOwc8s8pxQflWTMKeajhphduu9Bg8KCah+aF84CZoVC2Mcx7GXa4Bv5guaBol3HlP
Q+m1fmGRkAC9r/aLtVvDNaZuunse/VoHAcpWCpipQuWs02CDa5ewPVd+iMg+hlHMy3UVNpDqptAc
u9fBnmuPzvdv0qt5jFNJqg/AYJxqsS5JK3yljNF40BFKr2AZnCCoJl7QsAGHzN2s49VRC9Y6Feh9
HvBjRXgUsFbYMTtw/r7ihmW9K5u5VgAx7Urr9kfO/a3XxRUJ/Y28KPWZtbPCM+S10S6ofGwqSV/h
yo81oKMlfPNl9ayyCosre6bn0ao77xBwjTNf/W7lJeXtbQSwqLj6XmiZ3ZAAJ6KmR7Q6b4CXeaCG
fZIwRqDA5KqtaTxX9QAMrz381RU4qKVEI6LGsJzG9GLyYwzvrt39oLItYLKAHOkX0bzI6kKfgRh+
5NjrUl++WM7GQlglrKBAwmDZma1Uvm+c5EQFT/I6z3gi4+oBVK8RSVRVkUcqQDiIxVWlQ0pxsHlt
02A46y6Regc5XKBwnLBnKQXPrWY1dICnN4qxlywsvBT0BTC+zWkGgcnII6kuqw2SEInXkeVv8Yfy
tgShneKlDckfGW4bnTv6fgjHhbRWHG0WiPSxY2KAUW04+CkuOc7zoyl/KRFX6aibEXxox7kXP4BD
YG1bLa2ZJKkStYBTNrHNMnyH9uJiJX6ySUH8L/GX3IvcTCY3hD7eDPyYN1AU1T1TiWVhbOLvbgYD
M9ZB+gtBDI6xjfM1tsuohQqPWwRqNp+2E28AvjWl9kA/5ELxrN5iSjZD0fe9RzSPnXvqH+3ePunr
UGqDzf7rcMneF4YnXADpfSxFdw7rln6IphLrdXDhaDAh+cd2yWCe3ek07PmaUb0kJ57ZHrhn6mD8
n7Pd0gKhC/pMp8ZNC7OfLwV5m2q1WFduzsEGDBfBrw28e1aSH6oHCnFo4w5Me59LbV5jfus7PP/z
wrgtQ2spQNhMudOmLMDy4Us+CjurWkXnINTI5GpjljYkQSZYjS5khXWMRkJQbZi4OXKs4EO+qRrb
FhcfqwUzkYiR2HsRNmvXi756vft7kGFjY7+05JBW+RkzJJV6jHCLMz6/DwEuDoOJxzcvzWyjQpr/
GWFVt32Jkt8ZW2uuHc/2pUQqIy8TqBkSTuWr020jgOgvyqKmF91Z3fqKtw4kE1PkqKYuGcvem9HO
ZdPEYoQ5Ahe05pF68FxR2ag4kZ8huYridNNcRfsdwO9wJgYyMb1cJIy2cfckJSngl8ju/dUjuhSg
QFcZZAA0W19ldPqvkb8ymkygkX1HffS48H/ZHtsQKPmwX90x/Pg9m6rAw1k7z9gwL8jVjR7XWRIR
NftppHaflpDvq8OaXnWijVwDzAEIf/ZnEHxY7k/CHZSvDzvyA9oAVBnXXAfFbayEla11qh0fumoE
uy7ovxzTgjOq999FSAWnKio878r8XoCb3AOqdYHFcAlKIb2BgsQwHkC/sS08u62o7ZtUyD2s6t0y
4Yk4lLdjf/Ef3LEdfaXavO7kmxuzR2TiyoOGlKY9p/aJm2MKtw9Jk3jXvJbivY3jKBaQGML3ucAD
8bspsXEzJ44jm5AAXv1yrBHWJwXAMlCgmNQRzmZxdM14ecat0fgdmrs2SUGuzUHzJ4dIhChenTFt
ldaTW4QOSxfvU4WMdHyOtmYDRRJoY0+rdT09FDYZWncrwj75n3KSm9kbDXX8RXIhBUQj2sRBlZaR
tLwcMeYKEVgfNG6dfdVumv5s0+Q3HZ9rVkFgl3yWQuDhUmzcxVE0pqxzWl6q3vfB6+vM7+uwsTAP
kmJqYi1oa+FZsJf8Ic7lm1dd3J3cUy/mbdTMNEGLLxw9BnoA+GAW3B6CclKfCmxbFT8/QsaTtlZl
OoYLD1LW41wk19HwGQzI8YUVSnzwEFA24WVqdao5C59lUl5untb1/skKr/RrbreePoGLFEskNc5Z
VdXKw4nbydw254dZQbbgWFo8kxbo26Lt1dTglytMuLzNDWVygADpWR6/W96T1upplO91fdJdBqiB
0Y/s7KJEziDMlKjiZrxse4Yh0Q19kAes2rbD+6mCcGFbraPawZsSPoXa/wehPZE5QeULIL2Nhpka
CiJOB71k8x45eaqYlPTNGkkh5qNtSM+2FXnV6q90yHY+qzFA4N+xSEEyegU+liRbplyaaC1+MJNw
mptdx/pwGMSv2O0Aa7mV6RZUoh0WYtbN15YOzUgFySLKbiKk3OQ1LHbzAeax9MjsF7dyj4QX8G9W
i4W8DfSMpkxf/fP5IMN1E1XIPZN8Sa+Ts9y6qNwtdBc9NO78E7m8tphJMFMc+KSGvQDKQl3Bu+1/
fw3srZoWGohHi0+p4iULbqZOyQjMMZX9XIIXf22RMUoTaFt3C2FaOKQFzdTgY+l6cr2FwuID1luM
k8Y4skxADkQCcckESjKGN+8kIuQpVx3xFEMc3FEFZX1ZAq5Bj0SrYt7pu0j5FIdPpy8K397dFLiX
wDPGfb4J8PDTC+rZ8furhicaTkrd/51THn3ZB4YG8gGtYKIlLExRgxfnsPiEhbjX1ggSYlcWwc4V
s5z18ml+O5qlnN0GQAcDRUcL1rnuOUAvn35fq9EVP3++f9nB1DnlbTnqmMIPnVxf6MW/fFbXdNKK
VAEBeRDvGXxN1cWufNsL9LyCsfaUUKJcllSEY0HWK0S+EMxxBinoTdzN+eciCR8drEhYH1g/rOAJ
c/13XPjQhJegCUiZCUXp7bogOoJfLxYLFEYM1IuIDvAzQwri6lBAGjgi3jQKW6VQYJrWrgnjPN+u
2EV6cwovuKkcfYd6k5Fj60vAAqFKAKeJzXxTq1hfrGMP2MlydRxNfyVuSSTh+I4SQHInO3eAbACX
HLm5oNlXxGNsREHtxzogNIqPUYK+I7ypJizvYVFCRRpm1h60Q1CV5gkNmn8vK8RCfyGrhLGfmHMA
hMC+gBVIHcoz8YhSlIM0nddLd/g0uM0lnxdzqHwEbdrpPEJByesoY9TzRv4UQusPhc9kDg/sUesa
3nJuBNQ0E/HurwVXHxj/U8qC80QAcBJqDVsmQMYbwfpNWmdrX9yUHLo8TUxtxnoA8yFCmauoZSTr
GNYXx3aeuz0kfjemQpS2UOpviSeqWqq4u7J3VlXpRiJBxT2vO3xxO1p3/bQ0ajh7lPc+vVJUuV7i
iYwNfw5JojlJuPcsYGa3bTdPeDVK8UXvDzqZ6YSoKGnrVmVHcrMNPngy4JpJlHVbsg8k2AR08bAj
ffFNC3eN1D9KlSGTH6xBY4ZAHGbcZ6mhZM/SycKWcstOAAu2sSXxuDZ49UkHi+UtUav83U3x+NwA
qAgpcpZCPXEXe7yLIkAW7Him4sfZNagLQ5NPr8SqVBFF5pzXi1VKmSfaFjeZo8dCgUDsB6KTlmLa
RmaGY3BwfUMwyj5fnUfgUt3r2Si32X82XTN+JHWRRtAHJ6x0sqn7WC9RrIZsYridSLIAB7EjjJtr
cI6DDhKVwY/orlkppnbeXk7vcX1aXNx1IJQIYlUjZ6kjVaNtdd3zwQNLeKiaqqpi/Ny9OrZxfmH0
sVU6p3NQUrCVO3U3VUoRZfCRql2inaYP2cFbp4l3nhWVrX+EtypyBEtet/SqLwUwAnYzxkcjsSJw
PalAWeOjRUKR6aOsRTquPPDZcioC8NCEwt9i3AqzfPiXba8ruLV7mV/XPabYWKSLYkFqia0vS6gS
5FkS2dqRTGm39o8vY6qWkrXzKPNZISyU7/c5Gj1Vz4XNofQwB1dGpDXHYB0HThXT2INGImOouucx
s8XyMzdmhgGz/qIxxXGTVMcMNmD6v85Vsqc98ar8sDA1PG/88hUurjt6OgddsVSob2LDrJSuA1e4
guBLCK/aOYTbGpHjLk6jstHoh9FEEynP+YIA3aTdtu4y2R7u0/MWYs0Rsy082quGrg5OxqajsPxw
535FPQ57rGu2uSSOLleTrUsRHUxw6gKyRLN3UY3I7GMRhrOd//i4vS+R2uvNyX3OSubkkhFP3viu
K8lM+70LWl1igp9q1AJMybE2SRqGBiEcrxO1pl4W0mnovBGiQxYSvksXl5Qv5yQi49cZtORhKwce
XXE6EdwPgcW4jaiEZ35yfLu6QTV1uPLI/z3HvJteg1Y8gMTWQAyKoIBcligC7qRwRO6vkBBflxlG
ZVuqR2xpkwlSMTOxZGnyonyocltBd2XJz+1GLIOUxIGacxabHvFDsaw0tvzxaTaTeGe2936Z9MmI
AdyKKqlGwsT9AcyuYeM16XcIO8MsqbYNz5Ts3JLSrkbZamHbkndW6B+eoBkvbTglVQyZCTypkrXr
4hbT+bj1kNvXbXLrxqGXl1Hg2tezIvi+XOIaVLrzwMIS2x9k3K/iCTssmUBwDQhFJ9hyH8vD2xR9
PAFjxpOuoaFjVgQFaHm4zLUwxnxK9JVDr1RYztDZZKSsUM3L9XkZZsY/hM62q+lbcmOtymJ+XOTF
xzoJvMPQ+i2oC6I7PsC2yU3l052KCnVL7jWgUYlXBiDWCPNanhXoskC4oGqEHeKQeQgFTA2JrtDq
X3ia6jEH0BnYUovmKeMUfd4LR3dFLfU4u1EpY0ALPh3GE8Cp2Zm85C8Bm0O2NzeV+UpcUxzV2BPb
qmQloRKKrDqluBY3yvNOFOgFyPQ9iVg/neChgboazitXZ3fb+zHJRi0J3wLnBk5KKhLktXJkUyDs
3EvHeG/shLIiyy4+Pf67XRt4mojPrETpMPy01GjmXH/9ZujSDzfhz+CSxm8udA+fIQqlmM8zvww/
NrActXWHoGrtZ6WgmTA0lJN/CEtsj8nj0VC814GUqUwXuHeAaYPXjIoIVNEBS8FU/tu/4lMXAIgo
P+q1uiHsBxkLhSKhv9WPwxoiN8REkJHB3x90vYLbL11vDe5brTGPtFJxx0IquBmm2YJiTNXaKWjq
7iKj8r7zg2SPTszNThUUczll2j1B0XoSdAMkE0OcDMpZzMW3BrZ0KxOi+D/xWLBA2QeZXYXyg1X0
ZB1VBkp3+Km6Lak+TSXJ9idsrTgsA5O3TmwkbGl948asyZ214gJ0LHIkkRSXIjCGmZLtPhgFl+2i
PzY1XkuVAcv6yxWbGbdLjhX5cBKnrQ4vCvWItDi9sdiQiPum36Hn2xc0Jc/2HCG2dJIRZZ9cOP4y
9PQF1GSbx0qxFyYaTwUNnbHtY9VTrIOm/nHey7JZ699nmPeIVUJ2Pv1hP4nGNlDhCbHIEJRSAegf
NVH/PwU3jy3Bq5b1wHVAQKH6b8PXjn+oQBXr1FTt2mOHpgpr7WRbI70L/741g/YCfxtpKgIeRoq9
72oD4TPl9mxCdCVrGQe/xbsO5zae7idi6iCSyjSf1jvTxkdL/0fFnidPNFoNw9LmazNEgrcEqLRO
Lwgxrp7Jel+tkUH55tXDiCsMCSYDsRqeSBxYmeX6Ak12W/xeLFZwCl/cdW9CEmj7mUbm3ppwKuy8
cwDlSWBjaTdzvP1pX51xUSIHgB8IWFiFaCpC8MmhfcqHo9F4Z0rE8U1kOtyUNJYsuYBOxYyA/0vH
pj7sdcoG31rqW484Ij2y0YzDfUNNNfuANKbjFEVnOzgmEHD0L2t1+VWE8yyjGTtP03+bSTAhD1M8
5lNd1e499YRExoLNS5hVTmAjR3ISbcxumtNPdg8oR/cto5gWdU4MboYEY/nc4Oj/dZuAuhrhpS/U
luezW/pn/8KWSgk+vsLequjeKNwIXEWhMxz01Sa00jHotZPF4T8V/BkAj7Op4dLUtn9jJIWt4ab+
syeoau4ozN/VFpweYDhyfROydg/M2jnH6iTn6iIv9CAcEoXzsG9eBbZ0Xnhv7XF5A5VZ9StgW4iE
hF63D/x7DcpQZfFqWZ8yNzMivy1yCSOb5m4HIrvMPsP/nA4pAa98cw+/DUqA93O0HUDMqAzy4YAC
jsDLYLfDtlX3qC/DHArGvTGre/UD+7rlbhRxaShB1070gQ2SihZdfYRZjTnwImYYFfBtl9Woji1x
29tUK0hRxTzInkIhoblWTwlMFYzEiEyW3zPmo5E0zE6yHTJpf4gJN2E9PEpHARCvbpCUotFj2L3u
8EFkByknUFvsx7DGVrxHu+aF4ZvHm1R6bRFHb1DPDwBr+KtoXhzaplp8pThNtiIgaoIB/nJ+KZXs
UNB8kPttP3cmlneQAFrBvgw8Ru9fE9Q0+Frnsyk398WWyk+rGbD80tvDGrUIFJOq3c4oFfnFeGN8
56TWVUoqkK2WkqHqvsuRWoOewjrBrOOjFOtiyQlyawOhn+xf9tdHjkntnXLgnNdHuIBru523xL5a
g4Wy+yz2CMFc+lK6/xYMh9whUW75IYukPP8c9q3GX5lb6cUlkXZKAGX3caAGGsh2OVqM0AMCBtV1
TYdOEbA3yPidP4tJZc7VOaNrRDVwXZDK+ZqwdfR0KTepLX2OA5Iq505Rz6lpoJCsxoGNVqAggAq1
ht3sWOeZ1IDFgxeE5Y4vDO6DBzXqDfUrm2NiZU6kQiImJI6wtcbZXXi/IbwEShLCXGOjtrBrb8/T
4ltUwup5L1hxLEun8pG06q0d/8MYHbixdmSgYlmIipKMWvV1Icpy98a+/2rjYZqfkHMnE8Pg9ZY+
mzDzZPbgUGd28Jogsop0ONSgikaBhyikTEzaAPi88nXR+2DxYdtRuUHxKWXXcsapJ/vyUmcvBc5f
JmTacdJ3ACsKturnh+bBycNJnnAzglkeu+pABgNNGifSNYRPfMjLIrLesGiFSkO7amtZcvDG6YT7
JDjfcXSN30HcXD+ru+bp1PW54mNmZaHbjsVCDvP+yksfUj3Eepltw86Cprzx6rhFp0JhSr0J+j2i
lF95eJ7qvD9J8VSidOkJc3lrGsRebTDkXkPi5xyJbgOpzo+Ody3e3EK1i12FlSwm1ymZ3s7G80T0
NROVjYAB9EGE6UfqLKmp7zMLC0MxFZCcos7eUzIXVu+F0/lsUHM3/eZvIlU91Ra5ztWHQudYEW6B
PoJW5phbOHUqA0kmkwd72XmGx7YB2mSNc4Ga5YAf/L0VVRjwtZP/FUB1CH8Ne5pEO+i9ce5FW48B
fEE52ncEd75NS4ufo8c4HXqvNpZ658k5rsvNgJ1dAEYn7E3kKWLqs1sEZUmO4DH3QlfKjnlL3uEm
sKOOLngHV6ca9uLiP1ItczBReQMZeWo7+rvzvhhaM8jOujKZ6sbdwqSRlVZ05DEeAHVFoALkQwlh
3gLDFxZj4x0c0oDHIU0+1GcXl43PQQ3t1UWJ7DMERSyr/MHJDEgZb5LYE5q24Jqj49UOXsAf8blx
6e61INQNz3PZ1Cs/pqvyT4DxbmjwYI+V2MwNLEIwletkkmzlda2NneZuhIaXxZl5x1+cJuVn1RgY
LJsZfGXuBGe3k7Gic9olyrQ0JPia984syU7TEIVJof0b/Vg143nlMIGXdwA5r/rb4vKw9ZZS4hjv
7yLUNrDdC2J0evPWpds+ZjfPuf6/39mDCotf7Fa3zm83j+YHnNvxL4jxE7Dv/bUcNZ64oju84oGv
UMAUWPyYkyXTOLJBdS8Qx2ZAjVh6Ze2D9qdNoNHpaVY9pXlluJeJ4I2uuzX6+z/d56/j7nFxYLPG
ufRf7KHfnfGD4Kk2L/KrnvGqwNsPTojUNqwvz4BqkC4xZjVkrIzkuON4uqkc0PncO0nv666lFPpx
ZB4B+O71nIw9saFka+nIYQsbZQtUFgWeqjOLsFx0QzMT9ZqEzMH1m9+6QPtryaa1jC5VNOWQYUmC
OJBxXSKuupUTyezSZLdiKOnOS6AU6wEz8H9JEuDZdo3V3pBDatpZyP8fUR7Cu13w8EMTTEjUpN/0
5XOiB098CjJJIscvIsiYkbM1PcPKbDkJSiK3VkdniKzcNyxtGOqPGVlWeny9AyNUimwTii7/DuFg
yw/wlao+jY863+AR7YudkfqFoxp0mLwANoEt8K4vn5MbBMfWyxBDWiz85+obYkhmBxquZEhnMB0j
zswX2dT/8kZCxjvsYQ9Yly1gNSzWGwX7HseFYdhD0enzzyD0/l4V1hty01h8mkqUQehFiSNvlbUT
i4ZVqiFG3Gf0BxsSPptu9JrJcWYJ/VRTYT4c4kmjeSHoc/ZYpdc3v5sYSqyFtQFtEXP6sbcVCyR8
636xRGeWitkGQo0kGLegGzgUxVy3m9+4uynQJoRNxyXQC3UO48Jv+XqdMPcWNDNXqyqL8sr6dRhH
6LY/9Rj5jDB3F0JLQunncEarSiSak7P6rodWKkyMW8IY87nb7WNadblzJOrxVARMgf2lNB67ZRsQ
GXlMtMoU1Gfr+h0fhXB8Hy0x21Dk7s/MBh8NRYGCzyOZQ9u99rty+sKIyGUDU+AtnvVDSHt+U3iO
r7gjXIbWbzVxqSWTDD2KwrikEm956J9XDZ6dpOBQ83IlpYbvefEHTAxmCGYUaXQMXUZ59Osr6Gxr
sN5uyb8u2+++GrrtbsRHnE13noD5gSu0gL5LkndmJpCm35bu3n0YsdTO3TzKWDuMGSvPwfILPlEY
qY81U+blx+j+rv5ujg/Sb574P2Kr3XHAtRqoBTK1sKKYC/1rs8Vi3u/lWk4cceJXEq/1snKbcq4h
/+Hy1+SN4daUyurMmRokfqIZMzSSO/mdUdk9eq8QId2i0R79SvRmy313ggExZynC+DuCmnv+2fZ2
O6jsshXZtjUQnkubk66OE32yQXrXfy8ju31M6emPEF+ClPqdyN5uqrpsacFjANSt31Lq5pkC2LBe
jHd2x/bHF3pdkkK+cCrYqKEYT0OWDnLqE7FhJOLmP67zJLv/95CPtZncl22hhjpbuqRT2Qb+PlNG
se50dE/YZnmGzpMyZQ23jeC3llOnv9tIqxTUvYTyxYnifGPcPzoFJu40R0VbDZ3FaYjb40DfWWZ7
x7lA9FSHNxhyHjmFKv9q5qjDTssQMtj7wvOXvmbGq0yp+vWcu6G6DuWD/OdeNfPEyWy1N1ZjPZLe
BuCoGN15cbiDntBRk6kDtn4X9uP23wvnw9TajP8sGeIrGuY32Q499/2xpXS23BZotlDgYwAXb89j
RYMzQqA6dLn5GKOzc1CE01qyEn6t6ucnXECVsQAZFBoEc6Ds0FV3R8xdLegMD3a5aLNDCBg2Rlbe
1s0rRO8dtEkqG5CJGL/Z9KkF5l5DhiMiCnbIHkwHxDx44uFtp3qZN0F0OrNyYz7Mj9t4ZZ1OnWFy
F+6tjuPBm6huyJLUVvPMgjjj4CMCDyv6+i4Z5X5tYPoJxkrVWNR/MpvyV/578/CaiqvZOOKuw/G7
twxMZWm7gQy9MmSkh6QR+TlMjXFM9YFwHq38grHhxU4B6hKJaYtRzl5mLPfrwVWbrvlMK15xFIoM
o2KzAisfFeZqysOA/KZLkBKermyK0WzWQRf3YF/TS8Wv7wshGbeLJmAadUGs+Yd4Cak1qG9KBZxH
Fvcprri1ORVPRXg4EZH/ASf2qf9yY0D+iOPNXCV+k5mw3oONRaVpCJ7wu6r5T8bDE0ondWDX39gv
+aneUvkmMo3cyQrJCayXDzaxldM6L7zOPI0EtiSL+WR5GGfSpZWBilx77CKp2I/kMgkpmnzQ/Mkv
LVv6fniHZKIpPvAA/4dnzmYklv2Is+hkxgvr/kRG1XXayY+89CG1H1bcflmJFd4zVrf8Z6zulPqJ
TIswgrk0H8kwglRDmTd8OtNR8QmxwGeFQ8Ymn2XHAGs2ucgbs3hb0GxtLiLXncIKZ9EM/mIE+2E8
vNuzomx2/ODfzxWgpWSJ8aReRVkY6ajjiItdI8lHFn8+EJ5v05z2yyApE1XvCpNyBZViYG5WUVZO
RGTKoypQCZcd718dvJG++copZzBEXjRzsNn+eiZ9Wynl09E5KNGmZ4Pw7XMenGMTtmFIijaX6zwp
ldK7itpkQSQ3lAS8X8EHcShMcQt8R3rYdNFnypWKsw4W6OLK1J1vfroRD3V/AtncNiFzNgkQUHZU
ISGlVjwsvQoaSgHQaMey6y3TicZx2PbFhK3Kyttyi2wlW9WRz6NeycRhrEm1ifXVlF1+sBS9YvzK
XNZ/c+bOhPJpF79VuOkWs5XDaMOGT0QW0GV9uvHZKtfmtfKcVSb/lLA8W449OhVDU5rhKBDV1FNX
yE1hwwe0KMgUqjF8pRroGHz1M1V6Bz/eEDVx+Mr8baKCncI3KyRTYiAuWeJzyAeuEkXVzSkcfvnd
VwEvm8n/tFlFoRbHBOW8YS5LN7CGTOSwTn41miah5EfSrqIpyw0v0xv7TBrO4ELou7zlW/aXm5zq
LsgY+npQgFfBSgT24DQGawh7ocy3J08ZrgfchAcbBgY6+RqOBovbmg3dgh8q1uxs4aCJEvXfyfCi
RQLon20VnpwkzhKwzGe4SneopK6jMT3C0SzojG2fo9as828iqiGKYKO1H97iHzEw1m5Wr1m9OfQ/
NNatrMaNlwbE0kQ0g7rfssUdeHHtAuiDcMxEaQkSiPq3wzmZlC0eu1FeQbrNFTpqVmeuu0hI6R9v
L/KPjVgDABzGx2cgAyEvTugY8WwYARYiRbBZpHhoi57jpGne24712af4/v6jHupvJsx6mXbrTjCX
5kwgDtfUAVK9symBpQYq0bn1wY7vBCoeqoUW4pAs7h27kCkgCppKatmSCXCgCp1SvBr2P5IEZ8lS
VdP15h4qD2vS9J9LvByiY5zojCej5h0cxtjr6cQPq4oeb74c3FKe6zklfXhbHmz/y3rs6W/dakxk
f8luDtWSpwX3bNiD8tRh08Dlh65bxiSuXy52o5G3T9mdYj8il7Q2nIsgZUPEesIpzlncDQtdukXa
eOhmInrdQAiR2+dkDKJy46maX2csi9Hb7ZXtM1KT3wN8c4ieEEi0iz9ifYkSNXz5mF96tyC8kGQN
UFwSbvLX/z0wawrZ9Ytc0RPPTUPRRkynSaRv1EsWUBBK74kkYwRVOe3zWfErr/KwlVPfTX1OjgFV
GOETpT9gtHDJAvFLFHWAsynrhZe1mGSvBXunmgbIWMgnAdgK6T2Cx+K4AtltP0GJC4nR0uGiEI+K
51mWxZ6qdE+oX7LXpduFJK9TU0PVMdO7C+5S1jFn8QQbMepURZq8yk7+m72A2KihEsBw9KyWw1c8
FwuG+xBg7pQjZ+2G0rIQpQ9ZuFb3n2ftMkhpfX5PqT1pEfE7ec+7Mnyt+d2JaEeZQS9WiPpEO3Tm
EouNPWv7psn+qmQ0jRLC/YWff1vHHdpEJ0EI7t0VCKbhoORWuwVOtmKp8VxmjiwTSP1tbUejpjTR
ZMQXKjR9j4OHYd/AMuDsUH2NTEDHAp76FFmZQa1csCnQYFmM9VEz6NtwbXmlKUoytv5d8210JxcZ
AVCbMUHP5Jp/jr6K4Qxuh7dCFxmpBJ4WBev3U6xLe00hO/m1hUSP4UhJQTOH6z4kAfmfVVLmaYoJ
ta1Dmw83qYSulOfzT9PvHlY8r5frbsphWS6Qzk29ZTTj7KtBAKSVRYX5bTicdWhsJGTo81pIZBhf
AeipyZP4Nhb83T/o1vZ/ltikRS91d9bQ2jS0ywJd/hSQxzTghEhO/oKv37gPNJ8UUaZwR2MEDCeE
6Oxz/J7GVTRxQdHWff+8Lwtcjgn7GKyQ+XQnxTNTLnJ0qH6WwBe9ZiNHyyQ2vFVmSKA4K/MYJ0Aw
/VdMDhJOyhL+T1otC+vzVhsr4Fv02TIKRQW56sqe3mioIhWOlwVrmoLXfq/Em8TVVsbzgBbSrLaC
Lbf0qwGJ0nswBQrCAegNf/y9QKMh+u+aSa9yil3q3zf7tWSKWxFcFdQbax787OUkOD+I1+LjBF8b
GWD0zG0KHl9AhKi8XSp2tsEnwDa0CMiFPmfQC6A2AvDmSg8L0M2QE88Mpb9ko+Ewn2xv0Qi3pWoW
GWjGlyAMTyDs2asqdsJhNaksUBot62ua5fU5Y2+2MDKiQY2SHngglxJz+LAQQldUTLVsLkImLQZI
eP1HuNoAXU17pV6jzzYuT+3KhccvwFNP5EFVgEdc2b9aZ4XDPI3QKtkM2sosSmIR6XlPyIpK7e9t
cOzObP0Av+EvZtWxB8AsbNX9ZdqM/k71xKjVyTM/6SiYWpApYJI2l12mgUbvEW1zZkFOACFMxcCq
rvtCiUDiVqTfGII0tNUFleHHGX3D3glUM3whMzDJmD8leCAO3IaPXwElWEuXNtXAEH8+eqfegMme
Cn+E00qhbjm2FVEK/OqUsEkWSidxBwnnk+LmTRoxEdhGKeGOSTDnr1IkxIGGL4kvYH/6UFRqQjwq
WIYuVIWBdzl0p+qgnCKb8MGu1p2xmCnM4LnE1GRiSnDcn2i/HUhk2KkOKw5kNHd58sAnb7KeK9lw
tTkaFjO2T9XLgo+0JwWlwM7IbC4wOz+CDOHQagTyYGKBcLgsfX0L5jq72L8XOMLPnhx0J1v0miTH
rOnCkanLUu64K1EkzVhN9E3l3UBaIYIfPngS+nASL4XW+yeqoYuhOxVKmBrptJly58r7zeKDBNOr
DmoC5LdeeBbGnSi53RE026sfmfptJQJBJDL5j5DFY3eVOjtz8Hxj7/NYgiTqISZFsVeBFOhsOsC3
qMy0yWxPBs8Z6FQvf/IcngDO0TlAU7EZsEdFokdPUdzWax5DfegT3wfstAvKxcVeSA97Fs8uLbnR
tuBwurrdXktMWYLghG0Mqscv6+UpEFY0TFp7MXkqOEX6ScgTTGxdFapZSCdVyatYfQDKWDOPaCSy
X9hq0nHKXENerNdPYzITRGcq4XSO6KdaKwCoFnPGhkK7tTsbWAgtjnCF3wxf9wwrkeCj+Exfl6nW
kq7ccIO9fRHdhXwJuZr49mAPMF01lrg+WAy/uVtaEAgq9KdgJGhCUuLbvDCX9u5tS7ITFnpuUpgK
EhsgDVAs+QXHQLK1kKKhDJsoxSfAMEqAbEzA3eevl4bEmFrT4B0ujDdB4yCBt7BwFJzl72sKP91V
KdaKwEmKYAibDzTG3flTnJFaNo7kD8ed5zlZ04D9QEIFu4lQqJqrULFRECZye2CWVHOqGqxWKaGC
RGvjrPfbgSvD8QN1uvSsnHxpnRZW4XjCcWNKGehp4lPmfaWpcZGweEtEWyltNMX2nPB5MKQytvh/
Fq6h1xe6iAfzdcEwrOZvq17cYxacw4iv5LEVKHiryp+ivfRfSPiCgosR2S/Z2ITz1unCx5GmlPFV
HM1Bg0hDLBHUgyR7va/3WTIl+JsLu/kOjZAaAul4jFE3FLELAfkpLkp2m2VNBTXRtW4L15AWEkZy
LcBCIJ0lxwGNnOuC+TEV5oQjXeZX6mgbzEuz7jsMkx5wOFwb77d0wxl1aiYidTIn2RagskCs3xi7
371Ywu3V9BKC214F1Vu0AkuoUMyo37rDN2q1IrpZUTvfa/C+BPlY/8ozRGx7QnhGwjPScc3QIASb
/TjrDkJSHjUmT1QgQFMw/OMmQ92C2p7u908CHXooOQ/m1NBHrx6rhSP8Hzyzm0ZeB20SfKv8RLWA
v0EteCPv6RIlPoqAK9+XnBlX/r+RjQdV2iNTMcp3roxXOT0ZE/T++klvIspdMH8lTI8dkOawgDEC
DLMUgsLBCZU/v26/CfhWf7rSi2Hqb50qFxbeAkv0ivSakQXO5lujty6C3Sq6tqrFYXqdWnbj9vm4
m4IoYADUaSF3UBoH9ssoF00YaZA+T7ZpDUdpoR2Hbc2Qx9NP/9zRyN705UoOBXTY8e3xmTmicnOn
+1v/jq4upI3oXC9IwBQ6Hu9NyJwNBuZVQTUHvTpNC0JjmrK5ATeupJgDjp6t88Ivu8hXnt9Vpy/h
VrcwzFNqakCmGuhFeRXbLg75CU03gPr25XufRPskn2zFC3mUUMC0pY3qfN7lWzrrl69uOqgftDTU
orEPo4VVy8959GXWxQr538GPJ/HKNVTJj6hB4zHudPSUFhkhzyCrhdSej8eysG+m9IGUTeKYbuOV
giaWddyL0Z0qvJw+oQnbCgLY9G8kCICYxIg1j038/ef1GP65o4RiGBhNsRAx4RRTqh2pJmoyr4E0
Kdi93HiJ94mbmHPgX/IDmT2Xwc4BTnHhfM7ygy07HS6l/McCWq0N9fL+NmsQCwZKVyuu2WxydQDO
m7pja5YyY4EpLJEzDSQaaB8/K6kIpebD11Rh6NlYjWyWHUc1uno4e0t0piKRdMqvn4EqZ8FIAluo
5xj9b8DAVFq0u0pEyjNottzVxcrWV70msL88u9WP9F/vYiv3ilnS2vg/8I3VmmIGZB8B2idmFRS8
9cVcYbktolP+v+eEL9pFpMYonecz3GVYqFc2YNf6aoB2AZU3FxNdvjloz5qXy5hGKS3KeLwQle71
Em0DuZUuidYbboHBfOqapd1IGncEFxGc49IaOsVeSQmYWPHNYR+24Tfe5H4L+N3Q1XzghqyxIeEj
76MUbXMLDag7sBIZGMcDFyrb6nYXKL0Sk3OEsKtqyL9g8/MgaL1vI2extbtJpaR2EIb6UfV1B1JM
/31m1dfgKqWn0YMRqJql9023DJF9djh8550OLaa1B2hrqdmPYODxMVx5LjIrLHXy8gVSRWk+tXFS
dCgRKonqzZ/t4apfpnIei77hnd5K3FSnhQslPdHCrCOX5RYg4yPrqUhCDc9JpptsmeGgFf7EqZ/K
fH/mDMh6zI0wmSBiBy2eP/myb/cLNEN1oJke9D5B8uS9S0MzBWH0FoVjQnhSWQsY6I8m2tsWlhE7
QG9H4mwRWoNpTaUJfXEUN2iZYGYHw5Y/yHycRfa4mco4scxneWpldOggV47i+Sx2D2EveDHLOpi0
MceKPkaDfLke6wtvdpAwre5WdG110Nk+KwvYzgjaPR+46KCh0K2pimGH3k8bu4wtIAI22ogzgueY
slwlCf5YcjFzX3pskfG+bcGCKPK8hz1dSWSYSIQX0RLTRGd/NHaP7NgTgrKeeZzvDal9YBEuuWXx
gBDdDi+PyGy7SR+RC185S30u+HEOxvb/tqdc/EKc8s6Lj7bX2uC9BjCxa/hpGGwac7FBzsnmutRq
Yaxo2t8Qii/XrFBBGIkRJrtwmNbdQpgqZOezvD5QVjkPnN4KyoTsm8AaM/eFObXDKA++ENzg6v+n
Ypdkw7PtIEo+ae2JLekS6uZA7sM3cbJtrDVges8B5qT/0aITSHVLl/SJQ6MwoXTtLBepeYjknV8f
84Jt1zQaOTmNd3e0irwSZpEw1LiOjrYKdFV7FFnQSh3Nqua92Cw5nefaj9hnulsmbGu2r7PntnoX
AIHmHnGuPPAe3lHbpvr6F2Xxi0C7+DDBTmyeFZLJsKm1qpdXfS/ywrUqHRjQXv5kAUcYm/Kqsgi/
NnDxoQ58MoZI6mIPLbYOglekztiPJuwhPhd3Fp4sHxu9mhObIQq2FDgEUSQvfHQxiRzhTMCo4v2E
vcgQHtJeFUY5G3RHXcphimarrC481YvrVF2MQwFpci9SxU79drjpd+ZhWrx47bf6QBmBXHHbr2Kj
EtN565A12gYeqLny0rr/xnhCkdNf69psRizBh0NdiP40rulhZhNmtx18U3zP85CzhF3Frtee0leW
8K+KgF/El381nFTq4vUoWEvmujF0KgpQ6kMYJo6VPDuooBqxfHR9vbbELtP/iaz6et/khQXslMtO
1i12u+giIVJwSsty4B9dQUdV/2XvPbpnOzGbL0H1mIHez/a1mZI0855FHZUXer6by+Ib0QUIrSkl
u5MyuQJgY2U3fpNM3u6UVpdcOoLrkyrgGrTa6QegTJ9enq9y4LVbj0+7WGadBHaP/ImUhl8SWSod
BV+XsB19/4RAxbc+mLweNwhi0b3VC5NHzF2goulCv/gpMPQR1VX9OypK10DcJHt+SGYsCkmI8Wa1
C4qyjKA093zakQuKYQVSXmqHRpkWjHKuBao4BxUvxP9V+Xcgv1yf7+t7bd9na4y5gwMVfkKmgB0b
cdXr5TqT0tgSycIbSO44zrYkvrBTcWtqR2NQ2Wh+09t2xZihhqjZKcU9/kLeMMuZ8sFYNCtlN0Y+
qxO1mFsST+bLiXaD/PxBjv/dW8k6EqcwN3t9rd1wPUy+yqMeZZtnHF7X27/D5523QvQ0WLfIcfXv
+cauM/Wu9UI2qve1pJhifsVBb4HQ7Z3PMi3QxhFNWI9HHtqX1SnOJYnpePQh8zq/etmGH9HKnL+E
mvJ4Skral8ks3TWswA5NZ7LFoLBjvxx2I4rRVPzYxq1EV5cOGVFp5DKTepLPQQs0jK8FqVd3Mxnz
x36vdA638hicF+8PG6/F5yEcYexgvC3Mhec89RjOSouKP+w2T8XODGSNwXR1Nd9i/RjSQzpe0PBM
9ZexYde4bj0FRMyTTM9KpyrU7U7NOPFsCnnseY3ljP3zsXOTo+4hEoU/H0LNu60kRZZazmjeUpnO
sWAUjGVzm5rjtAoHx6gvKDZsrEu3A4C+rW03syxFrxSE4CB2AxcQH8OPeq7cZUuPp7XvoeVNbqyW
LO6sYXhoO704REvyT4N98p/LEhEKBYkQknmGzlBSkQLlUIx8txLSQRqLLz80zva4lx5HhIRfnJhs
qjo9Iy+k2T5vnQJ1bDrrqDhYpwqZYodLDkhkNiZb2VvkwDKz0XSJOAF9XxovWmRW4SRT7Ofkkd+e
bZa9+9+BCspqsRdHRW8v76vcwBKeQ/c0lzn+lO6NsSziRPk/8SR4CCHNrFd8F1WivMLm4Do4P8wq
dk1ekrWwBHxUU//NXYDIMXVnM6q3u55lzQdalsbWkCnrgtqD8aMQLrKVXuwaOdOtS/NXksINNOqI
S2+P0kIPnTCGhxl+2jYv6rsZUQ5XorHTDI3pJHTAkpOqvSaIZowv3++uOQYzMxhCQ1oi1/QJbHEZ
iX/Or9FyBWSj90qk8DQH8yuv1NLOPEi4D5hNitGfev3+eT+wpWBUPlxV3FTh30gJbABBEYeF6+Cj
FVZer4FMuhSERG9py45unP43S5kNswHZTPw2qrpPQrSYdJ6U+ma+cr6YmV+sX+UubfS1JECbW2Tj
7WlS86HZPgI8Th3GWlI3cNtwtFauwGA7SR9ElUSsGEW2peQy0biLP0htV9ll53AhDKSx3uqrB+hN
koLLJqMcy7g6ulyTCwOSY+x+u66h3hG1r9c4R16WL1Fe4VwLA/7kg8IIn0yjLDONy/NW8CzeoGlW
8ZE0cyNy01pCfTinVGdlbjhw+OCbhtEoEY89tW+CeTL/UZzNccRfDW8RBNF0vD+TDcTZ0UtjgkB6
O8CC4rdxefqrO0uSclbd9VKoY76UwKgdzexDNe3+8fSKa0l+ujVFerJwmAD5mhD1nrYPmdS0uD/P
k62/MraZhopHwaOSx3EbmLWJ/KLnnGisG1Bcx5j3kLHK8tCGNbYHJ0R/5b3LeGK688rwYwr9YUu1
3ce9SmVrkBsqQx0WbfFBYCZTwvA4TztETRRyRZqykQHC3tzIiWTF4hmUfeMTldCEkms24P4YZJ/x
+AQ+xMD2ISzQMpNjq20afSrXMN4LLZJa7gBhyiY1oEuxyxsVWFNWknUQPOzCjuTValPNl3DCGya3
InbTMzgG/e1Nib1YfWaFM0DZ3gZQoNzLlJ1ve2kVJw+lHYO6z2RsIUIFRnE3/ySIPgNHpfmUoj15
Udpt3bpDZnDu1Qci4hl3SVN5L7/019CZwAi88NRTkKV6Jj5r5fJokYT65ZfmsylsjJXtRFDJsVBL
GgquDtvXujPsPXB6PW3G8tYLR788cFX2gOylTE0yVkElGx83V7WM5wFdqN4MdHOUSvEFIta35dya
QEYGnOonZud3A9oG2OOsOB2mzqM5jwJWGDjljlTw8eSBuo4zazjU48lr0mt1K7O55kGtmaBwJGyj
iZtUa0O9YutWOLxt8GR1BYSoYlN8T7HaITu8/X24v1hRxWQrAmi94h/b9MP+d9U4Ah8NZhZmxhgF
Tdpbp4jPpwx9ZJseupwTxXkvuydhI48qiR00sHmSkzghCQp1v4nKf2ZVcSdR65SfwHfLtqn0FVNC
6p3KxJGBXZzojUekFYoBFkWNzXvbYdQsBYyQs4debqUKiwZZ7xLwpqDkSj+0LQ9toupkVvQBoItP
nAq9pWsb3DEfIpvKg9vGyxxMSSeJgWCWYtRESkrOD5sDWVHIHwhEldIbBiWRYCk8mqkgdOP9QYq5
XWPuxrgYGSuO05Vr8KtOEgxFyTDTb18UYFaxgws9MTb13hyAYfO7UxTFDZEtd7lvSgjjqQ5SaIzN
zKnnA2Q6cUY/2OSdHTVxJo6KfXaMu8jAUQr/vS3Jl6g8YfYo3ANYySBis2SAR4cF8NNkW/TRFD8D
y5pCLfulq4Rkk+udpyepDl8utLE8eRlomHCd0Zn4txPMx7z2kbciR9apc8DPI2ksx5vTZ9xgHPk3
uyfF0aE0Cg9r2uARYhHQhTfZTuq5Dvq5DaS4JIZPYmJUC+krEnk6JndMg/ZzzA6/icQVldUNctNv
9A6ejR13UyjcR38G+CJBN84IlkpyKcHZ3RMlvIwULp3fIBMgyLlM46rz+VM3YGXaURnlW6eUD6YQ
QoE6mu0moxE65zcK0+L9iN258HZGF6I5KMoQ5in9n0F+THRiQYM/bB8dxsJ15/8Wat5TZVxUmIpu
jo3jCUWopfexAoWko+QhqSq+7rVdipnpQNh7g5EevbVgXKN1ma7ull62HVEZtzbDS4L8nG7uzVVC
NxEUetK0z20OM/Y3vwRYiR1YXYG3SKt9oDORPC+IM6b9/vwpSblH27rrbpjebGlRuaHTvlJKzOjq
DT/B6Bkmq+gZljt+AGSJAKxIV+MaF/z26jDOScal+3KVxlrftNC1eQHFELpvyyqHjMntrAzuYmBW
guYTwVZyb+RqonMcVD3u28jeNDzWDGF+oGvFsepsk7C6UTCzFJFW7+i/JbS2dD6HQ6Kczmu5pAnp
vQJDsrKT1DsUCYdT+1EAyXKzF87iTjr4ZyBo3PD9O5Msz5mOA60FSKoJclxt0yWTB8QDhUgglCPu
7c1XyUF92iEPuARYnHi22ZpF94wmw82fEHhL2asvtQ1RLaZf/isSQtM4eTgpaZyEt5//MLmYKiEF
/JKQmwXLOUmo9txFD7yLj/MkyTHwkR4avwGrLWhm2G4Vr/SV/ciuHqQfao4WMIAM8+iRb0Kq11UG
gUGioPssOP6pScxPoSYOHzqt5c8yuRzzNCeIgeJFdcyvHgwA5NDp4l+Yp9uYWwRiaWiTzpAVN71j
CSpNs5gmgwxDorBj8k42zQjR5cGdpA5K2CBTo4As9YFPEQ08K9TBOglqY/IWUGyvAnedISYiN9sm
Mi/JQThJjPwYJhiP6zirvmJBDl4ngctNZSULr5OdWMhHu1WfFb4RqLqTaQU9E7iUl4jT32RInYd8
r6nAnwD6RHEBmkdLIpQCqzHYctq5fzs9Qv+kmhEYdRymDM5Y/hF3BE7TVnsCtIwqvcAgw3yGMba4
zeYsX2hZIzVG0e6mqSA2FC3uKhRWumUyZz5oYmXpMEw0FLLDPXjlp9msZCTNcYj5kieMKb7t8e3t
7eUvFjfq3QBIL7kQ5TwWkMP/tCfkngeyOJ+lBD5ReSowU4q/cbUvPQKldqcj/6lq3ECvLKmY8ajZ
RNzgN9YUZXieyli63ZYPG08DSOAXq2yFNvgQg9ub1GqMZEUaRQfcDh58MvfSK5jT/O3rrg6kfbaj
KcPUUX5Epal1ADewQ1MrGBsEuWlcAThNSrsckjp81okVuVuNWqjc9D/wGKFGRBfhi7RUz8VTIz3l
hoFNm4xL13PY2ckrY1Maxja+sr4Srf2xN6DShQ7dzTovXdu9mgUdZ/p7cm7aVo39Kw9uZgqRCEBQ
8VnfcrE5m57CaZO5amRiuGQTqA4gyrbVng1bvjt1PfoG7RDzXKjJBmjMSSBuwByo8JOhqlw5dXc4
YNeliAEAA1bGI1+RwDGgD4SGAafGOtxN5cjTiMpC2iBhmsS/3sOPg7POFRNNkLwl9IqM6mjcztWv
nBo1h5Py6oE3O7Wi8XtBtCCgizhxK+UUtSpx1hKwTzWABJO+CY2yMyxt/ejuCb3uUXpeervFMEcD
f34S0DTVth51hfJcYBJPOfagR42LBVCOP9GkVCoGqDsdH3Y7BI0TKpxZQUoT6dHOkQJI7d8EVRlW
IFnw6dZstZ8/liRRH8h7qoRsrxafog0DKB4AVK8UtZggChzZuTHFYl9/nMGFk3+jMTBbl2Lx1SLy
/JzCFWDK4UZ8KnWIo+d41HksVcpTdqBNsN6P/ByeZvjAYrTip11118qsEoZr9mtaa5a3puHED7A/
8OdqIWKhy3fNWCXyMrPNN7esGbJc5wrJOuigZZti4CM0PMO2tgmhklmON1krJPpr1PvCpvnuNGiV
gASAh0NPPYoMJbvhJzl5252iA/vUfaF7TqB+7tlj6Xyd3/2R4eFwCeJ7PMOgiXNmJODjT6EftpiB
NUnKZ0tbf7oQt2B4V99+LwYG89qs5EIoGpBJCiuFz5RuxnCM0qeCl+pakmHLDsGKL01VMsnwJxvY
yVLaI2rOQb/LgzXg8P4dMCaP1YmxonG/9aaCMgTfxDmi5Ktm67fHWCr2ISD8vQZ1G0+ypiSapSsC
/MHUsR6h4ZIsfjYciZe1/68gSLpBZV6HCRXY7AgRlsX3EXVMTG9NEgthMypQdczImZ1/jxzuoIzG
hY/B6pSba2Cj/x2TO84UQu2iRTPUdvFNLVHJkGnvo3v61PMv/pBCN+FcfDd7YbFj6ktmXjXybHRK
gkoFak/D2xIDnTDHT2PTEi7mcxLzltjGnjPtwjakuJG/Q/vD2vEk0dE30uksNBbVEBuVHGDn3niK
RGN4xKVEbz8jEv/nzFucBEQ0sCoHmGi5Drf3agsbibV15TZasXLmCLvOZlVGNDPaOYdVAUVdSY6C
23YP6pgZfmTqbZ20nvwuqJeNjqJ6hCg/37H5hzYtzW+xasvk6BfGoVXGQNwnBMinK+BB21SxPfmX
g87WG4hYbInNEvtsq6GwdcKbDklkoK3fwLdEassihjxXu/hzOzniWJphgzDtpXGD5h67IvIizpdx
DS8JbERUnjasZmckbd6t9qEV9a2Edrl0ySq+23qxxcbjHeCpqWu2vPDl5iwZjETl63jq1xgwHk+H
wroOoNojg+t8d/0+FyGBvAwYE8ch6VMgqr+TULG+mSqTh6Ng2Zj3ab5d4zRz+t9Kd2EmZ+BwVf3p
lIJPsOhVC5Ap7yTKhOaZ8PJWz/znprqb2+zIlaNtaAvykxPWiK6keYimg8rvGJebul9+PNv5GfAr
B+fqaeOcvhViRWGQ1bSRuSYoES1+VhjiA4iyheuhxDoFv43zN4X+x3skleKT5QSlq/3PsKIbLNb8
BhIBojgr56ydloXdLnHQgtgJWGkWNvnkRRk1CLF7SKfxbQZepxQhpNK8jn4KO9/UrVp3dvDLksXl
GmnKLZmJQpIHdh6zXCSyMPQSFPibX9HI4/nP+ilC1/YXZYffpylGFtN2Em+1nrnpjH89o/Zp03O7
JA1xmfXYsX3LVX0AZHTCxwN719O3fA8Tayy+SiAlHDe2a/cu/4gHMpojgvj1wXFfLDnJze8IIjmA
J36MxFD939Z2Aql7oTf6GLwWKdJfFDW3WsJrMzcPTQLy2qgSml86BpKpYPCBl3u9NF4s/gxCE3Fr
DIjrZUpGw+C6b5hEQP7bWP4j4jeHMpNDzGo1Gn2YnLNVF1L7iXYTRukVSwlhx6ccpC+Nk+7KnvfU
wO261BxU5ydplnCoJjZoAabIEpoDQpuP7JkSt02RoUu4HshNLHEatOJP5SfzrED3ef7wxDeMIG8q
KpAjWLwjJ5Phvl2hBJ/Vx+5I9SkL5bdgbK+kdM9A34aJrcu/8ocyo5qZdk6gYkbi+v/ly0qzqIM2
yzFFMGLAMz1WMWB4IoRbimszfMp5z4QBC8Nrk0f1nzcOUFxa4fv2ZXRUjev2sEFpEMhzt1uOrn9T
Z+dpPc4c3yfY1bePUuUwBuDM09Gfk0/2yfll7l5vj5r22aAzA3qQ+gp8gUQYrl1k51ouET/pUqVj
O9jnG91YzByzgPsrwYGaZqs6PdBklPJWWMDOGN//DgiDaUduD9/8/4bEGe+ccel9nzn0FKZnQ6cU
g7qUPk0khsd3iFknW5+GypCGyva62Qdh3JWuz5XxHmLp9kZJqLNk0wtcIL8bNAvnrq1Hs8IxcbAJ
ayvoLq1TsQQMcHvHVWvjLAV0oFCRnP/OPDiOanocB85sfvLK71VFgjhJDcZvzxyfjnCghPQufSjC
01OG365k4Dpa9juUqrgBb6vV9MWySCHrScVpKYTZtSLCCb8oOoZ1ELvbj69hCrW2h2tABIx5qkI3
jE4GrYt9ugt1juOlDZt+Rt3iEw6fWSNfcC57E2qPYzGZcZQFZW7OYTsfFG0HW7Q+41sjdjOEibai
5bWmWgu7oZCRv5OOHiWHMSIdtwQWquX5C5x368z7bT3SxF17nD2k++G8OK6ZCnjcf3hKcX7Y+tOX
+18tdjfQGDXNV0mb9H8msC24zbM8d+W3zEg9OULgiL3j4UO3Q7bmKTKbiWKV8vhQBF2joFc6tLuf
lzeu9I4LL51fMM6yCRdMUm6NjKi7AHmMq+YUbZ5VhbYYExI910GsYxtp3V9GsrWVyfQE+8b+aEzO
mIJyiOLPaq5yh6z/S+VSZt5nhphqyfPmfn0f3JRA7nWon8Va04LkjFsN8GknR3OsULCvEOZkzHWB
tbn8Tq9YG0qMdFxDc41OET5pAKJdhYF2uUk3GNyq1AI6R9f7hFaSHj03Wkov1joSZQsRlwQB+4f4
DFKKEK9pzkNSzsnT3rLq1yVm8w+a4VpqhskR8iq1g8QcsIPfWHMA34REe2nuVIVSBTg9jSwPFMAC
o7Px7zh0NPcbRd/rfiWy8fPHkO5N0suW2Vcm8pymMDDMth1X84/fOi0s/NGyEXxSi86/J7nYJBOY
6L1WKF5/icD2CV74nq9LzikFWCAPHIqm7npGISj5yyKvBt0fdpEQ2ObBGRaRLuQG1ofEsOxBOq0s
npCBDMrJh2a9X6grJFgvys3aY/8QJlzDhKXkuK2R+Ii3wmyKOZIuk28qIImIxTsgnfZ7udqHvjAF
tUFpi1B8SIdKONPom7b0pkbZirkrov4t4ZDL8o+NA7GF/aP5SV9RQqEbSSfcv4hzQQ8UD3zNfm3c
xy9OXeZ9CRo/SxcCWsWE/aMBAxazXlM4ryE8p9tSyu7WRiviRoGUgze74VmraJwRa8e2JFC0FNUZ
bdahrC91ZnWkn/0z2mbSYl1xDvYUDVq6EFmh4UkMdjKSqlOTHSSlogPn/0ETdxa4yGFAQm+Xt0Qg
MXnDRwtpaOF+snANb5cF4bySX6ZqwXNrOPfkwsgqDCBrsgBzjTcTcyfkb8yVYQVVfoI5egUqhA6h
5UTIWlZDhp6a+UU8/qmKt69MUxY0oTXNKUNYuyOIV2anjDXCJpCI+qbSLgRH5L1ksdVMwHbPfMYj
ZTHR+jjJGYAMGeSMs9Keg9I5KmLarNUzmqcHVVTBTVrZwW/888wmMxyf9aVVBjH8rOe39JvyGdE9
XTPMjTOGoos7HlxhqdZpU4mqcbQClNx1i6lLchUQ2Tlyuat0cAq1HiQ2JhHxiYUF6oRCRV5E7vHz
e1OcPHfQlJxe9i0h4evsUL7lNjZotLxSN5+EkdyFs94fGqiaBJxkXhm9XDpNLG08GclNRlucjKr3
tdh4PVRPvc24JOqo9aaUWi8LSliyiMLzWCCn2r06CeirQrHiYgdLS/FNb7Z7zx70Kq9q5r1u81q7
TVAGvvDPSfGjpdXu540O4elgaZ2CFSG2m6obUflDvgAK2fXYSkJKF1QBxqMFY7x5HYP3yzdLJ86m
EG5XU8v0LA8VJ1w6n7RXELo1IM4+MdvRbtKe+zIL42u2QbbHMZszsINmE4kU5ZbTJQXNDau135jB
Qx9vGMznRZKXSWw5pHI8kAhoR7Kn1JL28M0VFh4Mnkffm+FmX+WyrdEcdvf+k1jlzDDILnhnx6Y3
LAzxXGCcSU/ZiX+McUr7qvXlpGv4xj9++MiQmnmQMtPi6MCczaMkMrC7KldbXAXNorafdIilmqok
ZFYpVv9Fu0rQtc26/hLgnkj5HQPd9jV5IbYSdKKtsWJ5QR5BVrzPLR8xb+o4NcHX4gDsplkpMKN0
JwlfyZWXkj63c7V2oN4wfLNrP3/LPZlHjzfH8LpjBxDp7eJH+2PcoltPyrmH7MKl9ueaGSG4kLyf
a0/89znxYMC8Y7UcK0PHSAU/meWjc6dO//ecH8COUnGqsJDFunCFp2yANortI7dX0BlVYh/Ojp9o
+EfLnrqCyee9Osj1IHhY7cJ2tcorR/a3PA85VLDUL5n8uDvkwDkOo7gWVh7HbBANWe2lWwoZLiLd
6Q5mAafVV2HKc7spIcsV6KIL0zY4tuKsRiheK3DqXAWOlWyYKUFgg4W5H210uC79bA3kW0ELSZcG
1EnY95vCCzSsog+mR5L1F9dawEej/7twaGYS4Aiu/m03Njh4+OpB6brqD3D8z7YSdDSiDZuvmNjQ
7O0I55/06JDd5BOmusZrs4WDr7zLRTO0G3IOP88/D8RRNsC56CT/6wi0Dvt1sKzrRTIJKOIjmO57
R7t2n5/28gpmiK45kPzJ0wKYsm0c0w0vnRQC5OdDFeZdzBMUnAdR8feaqcaNeagwCzpGsVmEhsQQ
DxRtKvtYStPKwByQbYyBHJSEafTIojnClo0tD9VygRXDZYVtyAQ3upywcmqA+9/Sm1P9GzVy+uFp
+K87LjAoGD/RNoFjhIG1xv54I6+7OH7X7R0nlx9PWxQ44i6uZgBvQ1c+bCADIFLyBlJfoVEOOiGX
w9ovzoOkOHZKQXKx639WkqxCApJP8VhIjd7jhNQK9YU4M6zxFg6MTmpA89ZTYlhb8719ibL3mF2q
4eFAAM+feBnMVcDbiNZzAq7mlx6CKSBiGtpIuUyEVGrGKVPLZxXUzLu+f1c2dEFu4H6Ab5fDthgR
hnsAE8zgeQKQYE5CdNumvYKk3GYXmvKderOtPSa899Sjh/SVJ9d6HLAL1vjuzI7RHbp8uF0bfGIB
Dk0LYkuvABPezHdJqRDPKWav08tMySoadM5mF5weC5XVTELNhBqU9j0MaYFr1A9bP2qwKKM7JKdF
fr1ygpZvX5gMQnfaiM/XON179yyl/NQ1ktX49hO69PW6xR7+TV46sTJym0FukdtbP2BZRhSs48wm
+RXOmm3BiOLFf2npkhoGZ9G9ZLnmdiQvJMpfVb5uhoPgOFJJ/MyLuXnjFZR+DLqUQsOkjOo+uacN
eHByJYAKrWTtOPNlEk0KczJ1B+hmlnlzZhhjRJ5RRVzC2eYVcRQ5zNYi83n7DbS4MLg7KNmz3uOv
daxSLjGWjUcBqVQnDlVX59z4elyZORoWxaeBzWWcPpTw3o4K/o6Po64pvoe3iXt+H20yofEJO73o
1y0GzAIDwUdJ5eulbJXto8fVdl+fapsUol2G0TszCvGiIjatN6DbnDFRqENx4Tqw9O+81RpDwXfi
uzFiRIj7+EmMtMRQyt8qWiChVc3n+Wfmjz8a4iSNrQ3MIm+ZeBu5isJEyiTAd4bCkKBsnLkBNRJl
5/+d2Bm2MKJoYcvsLr6zqWxj0JGRda0vf6ZEvgboyPy65qNDntzZfJ6TYH1eqBOq4Nay781vP6Y9
KeXBD5azZbc4TS6wNalcvnHmO9EjWJBnrzB1ssI6ni+er/ZniONPMm2f/RRswQHqOIc6JK8R8b3y
GKUgVwCPyuQfDlv8glOEQ9p1rzryerSKAgOqdYIbUnorZvvVwfdcIknFe5uOaisXREDBb7rS+e0X
Gwjku8VrpgWCSqfD5dY8RXx/mXr805Cfcbgr5V3jPX8Q7U/YdYtyI5Nsa6CuTWkr69mauu5g6+ME
8cUtJ+3AS5a0vSNCusa+WZzCo2wZy8kKWaRoAbQgIPUyva/rVaQ9t0Ya2yon4zbS9C2qGd/xGmC8
+TXkrSgRL8n6eAxBlSJqvlPZ2Ft75svKoMtUB/11bWTWh0wLCTxAydt6w3kglDlXx4tuULEoKE+Z
bLtVE40jRKHNbkIraL18NV9lMOpZR0tZBmgAEPJ6VKNmVO/0boP9ABQNj36/9I53D1FZoJgsWAO2
lwV4SeJzzXikIK0qAXhVPisPuZFdangafSHUH8v8AG3xjHEAz4AXwMSXmYk09QqRxqIIze3MJAK0
i6pbE3KtOKF1l3iT3mL3JhBRLJYd81WJJJ6QaM/QG59uWRFY7scGiQjXkwdIjt+sScHLM9IqifFd
1hNthLPvAbbnHUNloT+ehn6AVPg0G8fmQs2kNiIbX41BRttiHlQeHCziLsH9NoikP3vKJ+xGOadk
CnTrFTI2NEM9R9PEnx55NR3Y559GxQ8raTlfXdkd9Y6vxT+zzT0hBxuCmkRWFrHDn7PdDvHIjyn5
x2QOZU1e3xaPdDd0ePdKHgpKt2yAjH9pR54A2r6VwRnmBm64kMixQfEjV0kyAkgnE2npuQR7pF87
GofRyvC5YMeA6gET+yZreUjgf/11zoFPXzmZyXF7VuSa5DJp9U1sVLEi2e64ErNHwmqSrUay9dk0
Ni5aDz/qc3yGejx5kLb3reF0Tt6zsOfKayU0gBGzjdBGlgRKVRyZEBXoxJSebVqXdMzqCJR1rUVf
C9fmZ3ZeMhmow7CI6FBcmrkojhTYxJuXDCVi28h17f9yo/AhSICaeBIi5ldSsC/36Or4lmwcLYgJ
Ih/rnLGPPt6533xjQ4VfjTNdlliUGGYLdQvzn/SKYxtd9rJu11QgVfNjhdueVMZPwUZ4QQQ6n0mm
FjoOegAj/Z4WpBegnQZegmY06kLTy9Ul1TKZra+EkO9MHArjSzcekN+jTm7Gv+IPDwwfo72TWBkV
T14Wq/bcjcEZfF31T/ERllZ5wFpDCiRXOlQE8GTM0IR4cCzSBpk4oGAEtTtw6saAUtEwq2ABSyZW
+jqOft7dB4mdhfEY/l3xdWURntQDpFLJ7yd92qSOVLeXmXTyPaVARUiPC58X+TySjJkwXzfT+sDc
jWYh6Pmj+v3kJyIIBkHboWS5lze78FtBsM12QJ4KKjud1tRb8YqtL+442ruAxG7kEGcbcWxZHU3H
u7GdDIRTdtEm7GWPIV4pXZXdPBsB668mN+OElkAPWb373qwqfMSLYSg1UD5W0rGNL/BbCdJiqkwV
Yl5wEPU/wHjwLRQrV+x5N+FjfNzBsGoACpciwxfJl9EMsj8I9qZIbg2ooc1NvSHLxdjH5S4VEQTu
BZVgRGorfgylPSvJ8EWyMud1M7lUbA4NLvNPxd48qLQO/YnjXkLn2etXpghUYtiP24OyE2Agx7i7
Dj1QCE3AoqKp18dsSLP8ZiVB/VuFXIfHM0C477YQqs3LmcXwALKYFv2qLmayQSi1jmy0DLXwdb1T
T6vna53ykX9Re0c2JSer0EBKLR6dsByCcO9ptouNjQnW49edwYe4glqx1qufHbQr+OTb3fm+eDLC
Ye4e2NPpt5/7Hsp/d5a/0QJRvl5UFdVQEFO4v8yIZIEY/MrY2Zf0Yu1CzoTtcgvDhDDe0yJvDWWs
ZJX7m6PKXCl6L6JvciQiolH0RmDc7hpMM6FUt5My5yLWtRRnvM86EhyD7g0P9nB12n/9c1Yy+V+A
UdNn8x+K7cvFY0NCFkULGSGLkyGf4xqoC9u+KdywoT/sPnwNqSyk8jbwmCdAFpHWrugXJDBdagGR
vlMHsJgVWmhQwJid4n3M0QOzwHkZ3Z3SpkVqsjO6Q43Dmvrn5Cjbuq7pgWtDnwM6UYOVQkUe0yDq
VstLMWtmqwsqIWaVby5xS/CKb8ZSH76mcmZeO8O+yyCZKEtDEwAj9XMf9cZqe6rMKmqguJ99fCHX
08hHx9iw2pEO9LZmKCOcmAxfxYcFKNPbUvQyAhu827HXMTM7hgT5gKYIHyaIzlqZW/CHxPiNOugR
dCE6OFbM1dXsFQdvrPXFWU+IyD2YFsCYZRSmRJd9O26q+2sKjbgX9hfxNA21+TrlX74x8nQ7K1Li
czCuhzqv4l85a0v4Bx7spznUtKeYR9qkvfw3E1vJN5VS2YNn4Xy+VSS0eY/fMesEPO/lIWPpzVPV
/tCWpEcWipReKdqX/xMWTsGGcPGMQ4dwq1KIB6bq6QftK2oyHWdqjX+enD4lRSZA6AuZx9yW5IdK
vsXpbwxjybWilcu7j/5gd1Z/s37j7k5CsfuHbqC9syUK15rUPIuxA/1EVG7HtAzE5dkaM/+IBVUG
7ArcAPEM+0q4IXJUjM5OKhvTvWA9lgVc2e2ItR4ZR8BPB+nfGMZAz4BD50ze7aC19en5iq+ETpsn
SMEatTYle8rgCv746uDg8ABpX7gMkcGTvPRxrM0s7ONwUv5haLwbxxr2a3ww0nUsxPmFOWb7VADg
V9H758qVq43FYvhGUQekzb1SGnFKOAhF2vH3JT2cEcWNL2mphRGGUzDUu6dzNdM3r0QztAVpC6E4
8z+bZQopQepjYV5AhsgUgvLJiyIujscDHFIwb4KrFDGyBB7A+CmRT3Ih2JgZTE4vn/ZICUYnlqbK
8zMv1z/Zcr8zQY2MHWBt0VSTyzm28MFQl6KpWDVr2LJBE0v+h4XJq/MPvOi/CASFa0WI8jWKsy51
lyJwtt+5EeG5YQosCO26+hF/vtjtqFRYXCXnvrkDSSjJkRufvFbAfV1Q5EUq8IBN5UR/gb+NgqoL
ET2Loa/IuLxOWWoh+Jd5YIBvBEJBEaCNECtTHYs8kFdPXZ23Mworv4QJFrpM1TXlHk80+/1tORjs
TuHxVbseJ2yO17HUCbl24wSO+hxUyDJpKrqD2DS/ScV3IWuf/ktL1NEFRuDhy58P50GI7so+v/OX
ijEggpqf6tDnLmGLVCyLQCGHCZUKn+1UH7PzNCUH+I8ILFG20qBu2wAb6H87axo/6RsxNqGeuQWl
i++Gux1qEcekReV/i2Ds9Xh20NDAM2MNb5o5x0g6equ08+rctuOWCRh3/wuq5SXx0Sw0GNFcUk80
lgZXHvixLvOfyZksKfu9UUwDv0sHhReCphz4WY6oQkDvQ08kderZ46OZDbN8LTBLm2ZzYh0O0tSd
BypjrTIGWdBaHihe+GSk07dlHqzExctRRmq5xXF10nE853m3sLPEzordhIkqfxJfr93pXJc3dMUk
MiyfKFK0IqYIOkGbwbiPPdClgD9bpArEIouj8SgxnuoNZuff6jjYXT+K1tioMOYq1KnPPlWhLcH5
cA5j5GW5LAjaXG70WqSvHHr3gKdXSZCMPqFsw3S5F8z/zCI/KJ/ms+q2K6cN7IlobBjcGyp/fJP7
iMqVJgbEqFOU20gJohH5VZTNQoiFeuHYE/r4QdRpKv5TAx+Eygdvm5MziL5cQZzD1indB5CXwwOi
dQzM0r/EFiI3Uh1TQNydyKFoM3rZ4mGQXaQDVbS59TbHPQTu8ss9jiNYPpZ4Tf8cXz6BsNYlivuR
wdP3NT8i6ObwX1Dvv/ULdBsZwzm6ut8uhbxiE1xB7VHm2aFcFRWP5j2ShXGhG+ir10jbdUL7wecZ
n6dSCmya/wInSkgNN8WuxB9Bx1/HfpJagXsMjJfuaVH59hHKL3k2bNlTXoHhIednY7PZjRFcWhga
kbOIX+TZXfFKY645H9FgM9UKe67MwC6SKcSP3Fe4VLOuC6Cvyw80astPKjqtAa+ZcHELQbQbo4nA
iq/e0tONdoPbetWQSDV1SsJphwoKbzfew1N8FYGYhmZiP9kkc3l3Z5hV00Tg6LWEoBc5g5pinWd5
G88fXcBW2oaaBRgZFAQLatdxVeM0lmk5RlK4sN9b9N2vQurCxdEkLSapWmrL4tS3hJwwTiABWrYC
yJ91eE9eEpkugRG5Kdm3+nQiTI6c2xP+tPszmBxZtpqUh172XAQ6BYSKSiYNDcbi+jNl35sfOZHO
Fm4iB7qgpTpQt3F7iHenx3fTOlxkgEfEZbFCavkNE+1x5gjPkik0j+Vz4+Zbc7OqRlGF9GPMHfFw
1eUsF8zGc4ZPLAx1Stp+OD6cPSEctXfr03fm7cPiH9JdXcbws1+RuEqP9NAA0t1frDLCD+y443s1
sUUbyHdlrxiUpzGyFvKB7Ov5+KQBn1xBAfqp3cjJ4Zj1YbxCb84nambYp1k5JXTSQuNvcTZPDIsR
6MjRlUnUTSOqPIVHRFIsHeq7u5KcLLXymRyQao5o5c8WbfPI8+k6vM9FJNHtlG/y04v4Kjj264Mm
8vyIheZPyrjSs+4HW98hzb4gnWgSJf/1VyCweKkNStHFkNXOaFZcov+m1a+YMyYPDnHyrbrHcJRw
GncYBjm7kndwi9lTXSElepzvI0XwK74aJXtkeyPSVOvMWkd4KaQ21lwgOsD+Fr6p9klS+C15aDKW
ydBis6gf3AwehQSmhoMLIyf1CTNlHo6HTNAGz41rHWG0pDlyBp+ZB72OUP6aW7lSq2Shw9RwyUNN
eM8J61LqhbatqzHXF2Zv2jDncJFo0B0nZGjt2gyamWdNCupONxnidVHdGMNzV0kbQk2+KRbQuiEq
CrqyA/G9LCvLx3tkbbG0P/cOWZ9TIBRVy2kDo0/S/lif/Axelbb6WxeBllKdhXZQSaJfp4DViNgy
H1/ujFzwKMEizxv3LM8cxmEAuXCw9rIRquM6KUQh/leqrpbcT35pB6xqnmJXiMI5w4l8186yPJlo
bE21qR6KFzG6+yMrJGIW2zXUVu2gGt9+iuhaV5wPdfelNoWFv+STYYuaiYizFRrWl3bSz5aUsqJu
oMw46pQS1gbcSZ1cbGbRXFcdsW4WolkFgcPYEuSsrcmHd/0lG0+280WJLvascfKc40Y1fJdK3vBQ
cql4JQfGYb0k2lVIjyyIqVz/NYM909S93nd2UJAGrR5t6sqt0XW7f+AwWv9Odj3yuOgIl+GKvlrV
VMWEDyRx8NoNVonuaZgcKZBAkyJgkzh0+/yGOaxQCN1auRkLMee1zqHA3vCygcrk6sv9f/yMva6G
KrdJg/4Ua/wfiG8dziq+qHs+ifchHOTt3IscjtytUQpieeVn9L/vsK9oncs20M6ve1S47Zu+sYET
mWd1VpnhWGEKzlH7sdXXVfRw1pnXBmEXiRA4+1CAKdOLdbvDI0fQI2t7Rme0gwf1T4Vr6+uJ0voB
x0CFo4TJpG9VDlh6V3aLrE8U+9yoMNic3oEQB7cTfI+aURI1ezWbrwBXAXIZ+iY5E6OkCXQoF9BP
sge4k8p5OCZOqe8An7Vm8JUhO8y6j6f+BjyHI/WmwpICNxFz1qAJ8jPytXUDx+ktTpDM9DzGDHsr
DBb9jSbgUEJc6j7YFu9s01nMFb7Z6K4yhsit6KKkKMxf+gANDo7mxfWtk4IhQj6udqzRGd1JTAJg
4+yPqkcTL7RM28EtlXVjrxoGmgMgle6YnhNT4Pq/kuDkjymlYowZDRWPzcgX3LPWRUIcPDTWNdGi
t5UsOsCj8d+5UYyJPjgCMsVKqKGcKohYmiNUZfCLG7A7kcbWCon0hAXze90xWjFuMYYH0ZH8zJ3z
fEcbVvkAcwiTrbrVVMYnhKV1p8giLTkWHldcTrNtzj0NKYnbsOAEE003D3LJbgKNAepZF8jGGlyG
KPJksVtkjcEG2BlplacXX5QhzaLpDIv4qr6FDkHlZi9SYjlkZXXxOKh0Dq8d5aEGFNRc+cAAzlUX
RxIdnsVaTQOix4fnbBpq7/Dc+JoPSrWx3ktautX96E9R35LXlCh26LstkguXH/gzPChV3466fXi6
RWRSOBtKmaQk+sclQO7b21LCIpM6JUc961tqahyl3MoB0yLjpNqV9QyniNjm1VkP+KWUqsLEvW4h
aW7fVwzVy0M5NjFsx2NwxLrooYppDUHhp+Ribf3B4+OMaloWu6CyWhWnJdfDZTuHxU3bhH9nJC36
Z7W9MDao5B6tAdP6rN3p+W1SZBUFTJv4/X1GiDXinNbWk+kBksjvBprTd1Xs1AuXiNBPAJKj9Lal
YsiRxPOpkKlXmHJfjdfBPM+mKFhi3UqwqJITVZtjxy1swNXOUHmgqx0xYSrstBmtwYNv8ZYCasQt
T3k5PFLc9HI9fMEds3uoNzOJFsc69j8qHxn+bG6s3ZlzeJm6B0NcmLKy0wvsy2dWlZp7kGI3Ij7w
13IXVmC1F+/WBArSXaGZm/rW57XBmqTBvoQJ6hKZl72+j5gHyC/PFs0jL0kMyKYHJRoXD+AnYehg
UJKVd/GMLZ5LXLTk2ZF1uGfHu62T/zOAn1hbURYBBUQj9zpK/GOTB9x+oDBorCqNM4SaeYh/zhPC
La14IOiCYAyt16y2OEi7r9Bgb3WiwymN6e77E18HJDQkBojGf2xVe1mvkxkTasy7NoY3F2pVDA5n
VPALVlO6ebijJxQ123+Zol+6JMBnmrGhM/EKMryDZ+2M9mvorCnZCZHimedj7tb6cPo7koRzsmC4
xO2dfRltNdCVCVFiYUyxq9uV9OUNudclER0SZB973pjKb0nbNGAvRAdYmYS3VMg6bEgqRdeAtFNa
4qoawcIgvN4/8Q0RM2gmqUodfNg3P/ogBcWeTmmKbZayPUImItkqQmtg+vp8qG81OFl3GIJ9elsJ
R7y+kF0mVLshK8OB1m7/eFbLrp74DzqAESMDt+4gnQSr+L31PCY40aRkeXvSSWD6Ab6XNg9aRSD1
nyfDZ+Jh1ao7GAt11iATlkxgKUQjXQYg4/3lhBNK60VGRD5NhNBdQdUsoq3H9x8y6gHTmNSrPZ3E
VlqaiHVZb9RocjsoHvFiMFUC5La9i4Q6/NlsNZYKf5rEW11pBOsBeDQvQ9H0mrTz+r7qFGxjSlM6
HARlxtH135MrFEnvu1r1yiI1atBXXhpLmMk8MnrI1AoDY/v9pBfDPuxFSZe9LxYjmksha/7qvhDB
IapVmXxV8Q/6drJCj4WNOWH3rIZqQe+V5lUAYJyrzA4DaNnbgcPnGpyaxq+vdACTKhV9I+S7VAqd
RYoWthIv9IwxMdCAomz7wbpGxa8DFcGbZ+eOv1mobIUPNbDoRDQekrN6fpf5JELPqDoVgARybFQd
OSJU3ilvXKZgkVJ++q7Uh/lL8qgTE4HUbba7mRKYOOFeLWIdM5hnfPjPfgy5Xah9KqCLfkKAu+0/
a4tZSMtguAj9+49fVHZNgz/pnGkLWcwzv02ofmDkMiKZBaMq6MJBnMEByIs4j1SwIFhiLMby7Y9M
Pr44tnTJAnSkx8UjDP83oCjVhikWi5dHPRbUWHiSpoMYZITIRa5UJPb5xTekcQwH+md10PknhBY+
pj+qbDou6C2M5ro/qlNgiBpMUB7wUzQ02WPzSnG9ax8ShnDMj2T0xpESR84L3DgyMCRi5tvi+8bp
TebwRsMSCRZnrz+WjljuVDvjePaLXAMzGgl5gXMRu+VZ6gY5WmdGCQWroLX1qOeN8lAG34Y389kj
3dU+niiH+sUiBcToe6Ja80Cjsj9cXUOLfQS5DfTyoWArofm8cCn3XT/JBskemjr1dd3Hk3qvzCrF
Soi2p88wSCfMkp5bW3SM4ac6Y9sfS2wVtkGJvSVSAUQMbbbWiXv7HGnk9160bIUOMqCavc2FfSaq
/pN9bvfSsXHc/qEwwVvvFG7CkHxoDzv/mxuiaBhmcFTUAb7QuvkctFQ3Z4TAcMkX4h9iKlDwcY2F
NjuOSKJZRQJX+QbIopSKXMhp/dlRPeNTxxFXlTPdhErpZ8Cs1VPOeXBxLn+MtuzMH88YUVi091ct
lsEF7+71VDnhYFBv5GowYCii8Bj0nUwhMfYe9SPjbz9ApYzKfCsvyS/XSYhsPAOtrpz0s17uaHat
YjxC/3EsXAXNXZTdNaVMaCMrRlof3650ivLKnuiuSBTsDJi0RL9bKQ1Nbb9zyAAN7MGDFrjTeZ/d
meWviAcYoYrePlnfbKO16Lqj46zMZP6IBXVa8Lb9+aAzlTVsnROq0TsinTO+KeEPiRaBgahuyz7E
4lS7p7k792C9SrkRpq1IpMI/P8AzuGwLf+g4sqRSLAyyUsIMyGOb2cYx7iKpRR/bdm05WPEpOQV4
ViCmgs/fdzCez/elHinht4NB6hskgpmo0l9T7DdiDHuZzXOZ5Uop+cokxOH623ds5doIpvHayG+S
0qjVZRrI9CvSCuCrtqByzny6Uat7JgjpSqVVBbp7ddw2BOTFKcSysNrBelbOn9d0vA6agO/1e7an
CsWgwaLVA+8pcCsLVDf9ly6x4KYeQVS8skkaLkSOLplEfQ9FVr/QnPAO/Ii8C7KpiOaqnDkz1y0K
JWylb51joc039kl0815BqDXah9aDPTEzTcR6d/B/U9CC/YSpP0Hk1jpV++7v7vUAdecfnF//FQ3x
yMSgGYVWcA38G5uYZcFUJiovCksKNLEes47E0rgUjvtfcZqb0wokkLUH6a7pIfXv6FwTS18aKsRm
xZSHwdFX8+9fKoL4iWBhyrpY+d/IhsSI6orIQv8sHFGHkUf9QKeC26zcchX80AdYgwoaX36DHvyt
aoz2n6VqH97hSC5eHX5rBhvH6APpUI0xcM/m7MXPxw+Zq4LaMfoqsBXLYuFjBG193sCQq6Suiz+p
xr+oyPDukajYtKDFC1kzhrHY78tu0Sb4NOB0APh1vHLG+IALVASP47JT/y4GxyFDPN/hORJU8o2C
0sXkJbe/qHkK72cCYQWB3PjIw48qaBfibZLdjr8IpQYNtJxm27T2nEXIZZ5ZhrbIsi8hq0eq+T8k
q2t0WItxe6Jws7VbKBB1oER5iUwLvqJJfqPmeGn7CYP4vYotk075p4+BAO97xP/bkKHr9Csr7e3V
Tf5ETVwKSUXy5bIbY+3Kwn4MW67SUCDU72rhJl8osCtqt14iz4BIp8nELUt34l4/N8Ilg3ZJxtvp
PkFV4RpcPy5HxBabLoMRxuuOEFz8fevAxhf2a47KlDfcRqV7srbIzDRO+vYncGniJpfM5vK1+j5s
9J5WKvLalhfpvAIt5rlC+Fbc32ChO3Aqi3Kxp8w6K0G/oi4gpf2IAlZb36D113H+LzPb35nRG5MU
GPuTpLa+wqC8HvvJKbgZ2sbVySdraoUM9DVFpJZaS3jHj5H0jtfgg4apHTlQ4nGpD+StuLJvs5Uk
0q0mu2ynfdn9EZ/mjA9MLpAD+fFQMgV0lYeYOa4yVSDWLdZpxfWt4mfI2HwwGLPAPkFsnSpmcDs+
GjlVe9Q01p7HclsMvxD3UWfokAKJS47mUC45DvCSBz7IAu3Js/Sz4S8rLxd09xqlIx8jZDPpH9eS
x3i/s/VA39ni/w2IZF73XenT83zpsc8dvUzNxbAoxLh5F6IpK/tf7L/GtIhsNDZCUpM7Eoi+i1xi
lC96yKXO1AVbUuDV1StfsdZNX2DObGVwYmNmZeo0WGgFSXvFZAtTF86S858iS+sw7wP1nsmmOYrY
0zhmFUoijhuN78aBjXZ+lRLusNLub9mPIoGMWGBEvpzKfB8CKZffwT4/fioK1pQAbrFRe+YUqd/Y
huGhmKbBHBvthoSY06JuulCqHBocaaEgNPeDYcVKlTtqvQ0zPg3XM0EzU5KKHuSaTTRZWi/r0t9K
FmgXKjin8n1LadGbc2JpEflnE6SEIzhrpRSdjEI5Bl2j9RfFjkBNKWKtHu2HOFpRc4DvQRVRrKjL
HHmeWZkji9gKTI292iJ6kDeVGhgpbEAGiWKuGJvJMes+UK8AYfCLMDN5XgRxn7ih8GRh8y0Br0jJ
4L41XXKFRRBon5dAOLZI46WZeKB8dqxZEFc/B7rMc5H4b5lJYRXcaPnSSrY1gIjm2iZnFwb3cv6B
gc+JP3G/16jkE6jqLPaACb3JCElz7bNP466EEP1VC2dSjd6D3stxvT2rzdxtusMc35vJGDOkMDf8
54J1dQlPhCxaBGC+mtJVi4lHmxtmbt5p10PGFK0nmWRsa6tW/Klb/TE8uxDFD5fxr1TYy3dY7oqc
1X+XHJOjvMxM9/YC+jSpI/9d3gNgcZLi9TBb2jVmlZMvg9aRZkOxA9AtLDLo1M72Qv8krbb1q+UI
/69kRToFCOACV2rcBRAN7py9ayYydsLu68efMFEQDm/0nnU+YLejauZn9PUhobG7gCPY70sRPjxa
s0CwmZ25OY8CGlbSXUfZUVWisO+U8tdoKMpI1WY+z57u0AVFsv7Vy/Ao46jz/ZDQ+FVaBYRg6+yV
0JOXj2aUvqXnlvfjaue93c0QVzodkUAHCWXHlLtB/oK5wjsfSV2h+22XUmgdCWspCJkFXVNzdCx5
xFXhshJ2nzwes0+eYlOc0VvHWiYMOEFIiDmOZui5pfNMWONaWz3+yod8Kxx2wBKg1uiaFGgje7YH
u5pBMJ3/s0i2vgWzae2hpeBFtCDhbCeqRAGtdmxnMz4D6kSi/N5lDvpoClt2GUlJxU3Rw0DTffdz
UQyMOmlVq4YmHVHDUP2eOc/q4NPyBaOXY2Ia6PF9elw5nzy/m4zb9DbNkVCt3Qbz9b8sFSmQjmEy
83EykNK2mZ3JBfobGeIbgSGuexhMAlw/17S/gCVDystAY7quN8WJx4UQgrO9+AVBdOmliqu8/uSO
ePs/5QZ+kpl6poFGmXB3na4WGFcL8GHZoWSv4Nvfp9q3sweIah5ySTpM2kBs1Y0AgfqmNdR8Zq7d
O+PSMz0NXoQghy2NIdRLjIFHPoTitiGbSINFrQSSNRTJEwnmwycPP8hvi5DH7u/0tVgAD/UX5Pb7
mJPfN6wASfkR1SaFJX3nbob56l7rUFsCwfIc4kNJCRNgJCA+DNEHlGZ0yjF0eDmrGLULHv6KM1Fg
UK7BRqLFwZX597yoR9h4gzQwG2nb9BNgU4f/FihpqmsXDDul8JmLXnOsaohmfP2CH0Yt8woSZzZR
NabsJLuMLIlRywkB5pqw9cYoQkVgR+DGRsdlyrHWpyNnT7Krb0D1VLLPlE6pG5L1qISmwwXybkwZ
5w0f941TEIUjeFlVgfAgzTLR+mNyBJXzBy4YNNmbAl6m7eVGuk3++pcdqEGHHy1lXfX/JaoobcZc
zPRMH7lm9XloMd3Qy2YbtSVSQtrMNHK3r5F/w4Us0zTgUHzB1o2JtHzWomHQ3yiCIqsVVpyUpe6k
mj0gl3d8N0oU29+kziEdLthy7elc6KBZpcFU/RZhcfxCkiTf/yiRLaGHOqOKzoB76zB9rkRt7JmZ
Rv3MV4LDTjPDYnZcywMkt6T68RQWWN0vv6RkLubvB9dDmmvXC5DK7MpTDJ9f9Li0IJ5Ukv3vZtrp
3mm6TzVgyi+hQJ5JWONjUqIJlUXRA1mOUbp5l6evRfeIfhm4c5FPsYdSn0vzp5a9q/yD2BviGqrW
8Nw/pARaOMg1U+UBZI8909J18u1b7ltjKYsYBzwHcEA2SN+x2ajoWQqnGv99iL/AtsAkbcr2fmux
KaiR0TvetGHICY553G/1+oaKTgdtGlQ1Amx/MxuM1xhhgmSO3G9Al6O0fBeQXo8n4EjKf4FiXuFR
xEf/rCocdsSbp/mBAfYepj4r+Z3XbGZg3D0is+Nj+4FtlwU5G3U7UUo2IFfuQ7KayEMEe5Tv7sXT
e1xQhQZ4z0AoQ+Md1qTNpjrDeDCUpVxDO4BqCPWRkwdwPo0VwZY9iW1Xnz7th6prwpL4QMhREh6N
YtAbI3Wen9FZMgYJP1PWFyZULCF2g8q8fiwN7e5KvKusT0HLV9VXZac/2NZnN6162UXGXRIM7Xgc
Oh01PBi5TiP91gApCedPZKLftkekX9fju/QKvTUnf5h5LfZtFd2hM3eKEnZdVbdhQ+3toJf3aDtp
cKmf0WINNY5rhWgnxTidDVZZ8mSZ/Me12fLaj3OSAVZ0Dl/7MIumZamtNvtcWZMqkm9/dtyQoH6u
8ZbYK5/RsXey/yvwiEoJv/E7fSV4qTUG8p77jBrUum7oH3YDUEIemiEE0pVH9I+PmQfwsp88vHR6
AVVs6PtHGTHi1G87915m6gZSY7hNk3fLt9igsJWZ2vn0yLDTFdm85CxoTjZ3SKztRQYqtbDMm+DH
idpnai2Q9drebrbD/uRx/CeGE9CVjVMy65Wc6JVm3fLF4xuZtULx3IXCyLr6s74gXJyhfsp+UXEA
zSE7AF2kXs0ZExUez8mj1WhseT4VnK6t4FQ83weHxH0OiNdPT4d3NYsDtv9FaU8DJsN3FfUEdiG6
+C5V7T+UjZ1H+0M9qP9/l2Fpu7QhQstaeEGp4qM90keHMDP4mQxpNHs9d+G9vDd0/3ZVIkQtkunE
nE0jBle+SbawYSjlIkmt7SKRQQpkp6AD6Vw25evm6B+QSkvbWP0TCr8UHfyoBynEcCEjDyQLjkhe
FZpAv1W4Q/gJDAz8dsJF/7RS52GFKHq1sxG6dV7M0aydOYcsFenAUKWjVd4wgg2ZP+RzpSH51zi4
uQxz8K+jY3IV/3dBULWTyQkuGSup+tKyHDpvGW9ha0Lg0STjaW5gJybKwy68l8eSxTPpE6MhofQJ
faiGCgcvAR0ybYsi6lN2qARk1bPxjtKrTEtTs9WEbIfKlZ0lGhXBhT/36Y7RMxhnHUtlCMP+DRrx
K8+j7bK0wsf+/4ETKiveWxvq1AlXkxZGDqQgdNUN4CNYoHGr5pS1bbox3P7em23oxrD1SqD1JuOE
lM9DoQ4ncs19xErYdrWg+bP3Ihpd0MeTgurmzy7BmRdUCTiy9lcmxYLWXZEWsEOJJvcYd7arrIL/
ql1vnEzlOrS+ZZFhzAitfzMCxOw9W48URCTE/KvgiYpEFORS9Ycrh/+439YiNQD43hsmLTw4OxEI
g+leESkb1PSKI71IP35qor1M16vdjP4Akj0/veVxzCt700lheP3uonwjSHKhXC7hVajD2qw/AZJN
F18BbAV8MV28LhqyvwPt/C+R8Yar8SBDs5NiohRkamG1Tmx3wr3PkDFqy1uwOKixAUOucI6UlS05
XXsef/6D6EhwUWRC5Hogxn62ySawH1C/+0c6bxNsONZXKY6zR5H0Hlkq+O65ZEohi7MLH5ldMHQk
Yznw+djODBOG2ZXVquU+Lb0hd6gM7pR2UYRyGQ9V8aq47fGm0rdsQw26A6JyM7Cy5EfKg/voZ0Ep
tJbcSVub+mj9x7UiaNvv7u0xnLiDmdm4YEAI0/O5d5fnjTTLwDah/A4J6p1f9ic31m+gbIMF+Hqn
ngFXpEs6sbtUacL2uOSex6Fazljkyhj4XVKJmWJvhsiRbtJCz2rg2HYvfNh3Rf+nxgxs7bP6JkcB
OQSf829rIXMnDaaUqArx16k9uKtG7ZzbAwJS41zy0MzpBT5D3o7jFTKMeC42vkzcCLtlgwD+Z4Ft
w5aDwqWBBUL8uphaqz8lRsCKyYRxg2MXOi358F1CvG2oYyVXkzgazGlcKAVujZvGn6wupQhecvEv
HaQmE8xvsI7bKzmzlpbFxYsbTnpU0vS3qbtQHW4OfUu9Ycei/xIWAH8fcqJkuKywn/7iQc/TFWZR
88Y02ent/TQUMaKqA8//XgIC+Tp4aRGMXZl2bAwQw7rOyAoBI2o0pX1UPqfD2GapdYM4V2/qo7l5
tZ3hOW1EScsMG0mI6Q5+rV9pN9/W8X1tAnv7fUI7vM01YRh2LCKz4dx0tDdE1JtJLWSo3CsCCtrL
fg3DIzoNCd07RceouIR6rBfe78E6k+O3ni87j5EkHd5kL6VSUoq1iHFwRL8T/WFkltTXjpvk6/Y7
REBsXxrwJgiaxujt585GSkPgG6A4aQ/NY+KcEHvyw3Ai6ZNQcl+nczozajsmTNcD/qFLtLa8kHCl
3JRpMxTl35RXbWPkmia85vsviKlUmE3Fi1ZQ7Qsn7QBXcgdj4kDdCT8WPBkxkBuiyRcyiwFn4Gtj
er+962CKdSeOfQ5aMl+d5jhGCOowlCcaSh3qKHrGyirIKFRDvHOjX6c8H6uYhSTKnLjln0bO3NKU
yEjNsGiJcNEH28kujjtRhdV8v8ORlYmg76jxOALR1mKnNhF+YlFbi3qHhmWtV3TQtEGstfQXSWBN
pWy07xxREgcJrd19uVYEGh+SmKaatO/cphRnfFXPd5fQQThMKkQBX8Fde2OsIWNQH5zN8Ey56yUg
NjOtwPz6vtfFQVeuAUfyhxrR5tmFhN8BMfOPpCGCDmuqLQQGeCah9e9Tquz9hXPwL/d2FetPS2Xm
IxflxsVzRrwXRaVVLIf5xw0FLQpYAuPs0XbPFY7JqXw23jMp9tQvLa3U1oCQ8Bgmx9kQa1ORCRqj
/ls/LfDeZuOJLXfdWE+ZYJpvVPyXpMDhUstWdrZ5jnwP5gC8IFgTqcdIpbQuEjuPH3Vyfdm3qQOT
QlK1YcMVh0nwMT4nyHcw3O643buZg/OxKPVcVMHAMo84wnWoF3mnJNKM4/2nCcGkdPicg+GE+X+H
Gr4JmRPb66EyBih0StSKVIpZBh/3vjdiEP0ithTY6WZ7I/z+soE5VG2pspz577n3r4QlzvCsd9j7
Bosq8Z+JYhhMyK7xxJxBfM+TDzWzahdeaHAu0qpr6Oa67WBY3Z8BfxSgK1ORSE/cADDVaz71JrGu
puF4DMIPD1a38xI8ISzLAGKNBx+KCZMwhxQ+zlRoD5X5lSd1/E3aCr6mxZYgYH+7i8iH3cSEAnGp
TOZcNgh8UNGvwbcsnVWZcnZBtIABpo5e8zvCinl/A5BxFKUyLtS2hNYmad4+dHsdGuWgi5YlvVFQ
/gYeeqf7oP/yDcqVcIPjtHqssVg2/iX2X5ma2uMS1VIbJmt0/aUt+bqva5GTqDgKHifBmOaq1NJ4
ofEaziqbtyiH/xXcadZBQFmHETQrZUg//ZTDM625Ngzw7ysoIGihtlCReV/2oH3R8zmCpKgEf+Rt
/QbWpecc7XaApEtyR2QhxQhNTDykncSa5DzaaEiq0lO5MBVBBUB8DYekKRvNj8fADT8gDAUlh8lF
y78dOCyCxRrTlG3SP0YvYTav6wkeHOi0lw0bbn7LQ47Y1hwm4AY1ICKu7ry0T5ITFPGZHtBe13mN
SyBwuBt/6/UTuvJyLSt/JcxaVY3BkTa6iydJgh/2Cq6yPChbiQL/08MuQyLOWGcygX0IbrfvfGS/
HkOTfD1Fj1PZRmId78IHL1FdxSXsiRFKVwdEWnuAxP5YZ0NvSSSmnHY8DUfsk8X1k12ucfvOELAz
gwTmVi1xr2ZkGH39uNs1JtWL2TRrPTvbwuvOOt396CF6NKuqIhL+YSUKcuZ7hMj/D3hEeqgxc4Gw
xygOuWhA1eQHqiee2g6rwy2MN7SCn/Er8lJfnuGMSC5NTNY4WorTMju0AewQCIA/LkJeh/gH67p7
MWLtl+aQKbuQO70u57tfNpeHNwiDtQJajdIDViu873QUfNXk6T/sOtYdiqeOUvcbAdrjPslYWxOT
en8Wl1Ftfff/0AAaqbEGsQcKhwgawVcE3tLzsP3GE/quuGwm6YVgiaUcp99smwWL7GFcUieJ1SEB
ACR+7m10v7MUY+3iK2yEN7v/x9hSkuU3ccFTFv4zD91aH5it0Y2YHtSJ9wxt7B3cBCiQ71hoYAWF
xVvNMiQ59fRkwgHiwttpFGhRNMTe5IYy3uM+d/5DSEYUFnlQmwrE3Yx/I+GMWzHDwHJXoTa5yuOE
wKwdsUOo45dWuy2lO2bPeFS7nMUOcH92r4ibjy75xEX5iqD7MGt6FqKIdR95MAXY5b/YOrvyRbYZ
eTmLG6pkTVEFrbZJBFzG2wiK6R90MX4KUl4Tox4YkmAKY7X5Ajw3cF3iJavIyUj3Oz+aUMB8FakH
6qWP+b5Omns+MdOYAyfy5lgFCyI15sl3Q8xBj2b5fnzxDjxget3rvvltq6teUm/EFfISmPisn3Kz
VjmdmszAn1JeTSqgywKXJORiNkrecu7E+UI/+cOhMlIcpOfNC/tg/8/6E+3GDxbfZk9xqEANpgs5
60iKT1uXK6+d973RxAl3Ayab+dc0CoKhasosHWmbX682x5C+ovmdURaS4X3JnMGMZ/TJscvJTLbo
bdInzXliB6aCeuD8A/eRXJsPUs+NVIcq/4bJe6arswPNf+3MvSxMCh0ZSSjvZPmj47Oj5V4y/dJR
fqXpK3wzuyRReYN+E0g/Aqgpf74gQXtASSkjl+vQnmHHFr1AGtPHBYcPmGkjF8fcGZmes1oY3SFk
lHiW6Gzdksrdxv0MvtuioEljiyAoAySpTvcg/Yu+KjhfzEx7+/fN6Zgpr6KopPawAluox8fuoO+E
ZJ+Ay6OrS0vOAV2RHjvjlzWoH/cBlAQSUBGOPb+vOOqyw8vunGhGl0hUzs/44ocGHrI3hYhiqTFO
6SnbU4JKy/8yeZYdazv88vYFqng43WAxUjxiaZ9LbpdlK6uWOk1HuPKmOBJfNm+rUf8NWVliFI9S
rySj3lXtXzrEBSB2lnP4oc+H1nTzrazaT4sNpVhMSxCddnNTDrvHsS/wopKX+5WEe2f5XtF1LIgg
ajbI4Snlwyr5cJTUZkzBai1aj+6rexBGgLmC3d+tU7LRbixDnRWmW927Vo9cmv5qBFYYXWo8Qns+
/yUFeFuKToeNCtU9QdZncc+XIxJGN3oIRLVdwYplnj6tszm0G6xcTw+KcgtrWrdh1YEacEY1m/uM
ab/Pw86xIkFk5LBiqN3HjoNLH8slwdA/ucwWSCK1/aivDf2VyuOs4al4o8wuymmBOsP7yfwy8WGd
Rj5S9/gR2OcALxkl56dnXW0qLgBdhN/1bp02RTy5CuD+L1ign7GfjQRVX6uGAYZynzDCGwdEThuP
CTJ0StZat8C4p2ANPbOVG4oXp3fE8w8LrWTaqSyNkAGcuE17Kx2UMPpuGxgJaShsgTf8tTTWfsxi
w/HDgjbvbqNiascPVDbexMk21hC+sUYZ/CcufHZgd1vOasICO+XNnjVdEIKpJS9QuLgjFLqnNSZB
kTfXY69FYyaF4ocQwdCiC+gqpjHxc9bzKYqfcF/ndq9Z1XRLXJjcuaqfgRCaZP2IXmVXz+yxNxBi
aMlHCIWqmP6z7c9jMJaKrtbaT0e84KsTZ2YMSsagBDfd5LPtajj3FWUJKvYpneojv+Q4GuBzabQa
RqKe3+ZvVai9PWpr6nRAxt5xJKK9uKLlFM35h00vj3gwDcPVOydH7FsJeLCV+gT63QP8GRfuf35/
PfdnMWyLxHJfrPUv6Dazd+ul3oXwqenY2BhZ6gyLbIcq40EYrHBzvZdrlwkGULncFso0AyI5AHev
KWwDO5gXs/6KC5sgeRu86mQZfkE1pJhPTbHcKC3FGd5MpEYaMw9gScPN68Cf58IWxvhAQVkjaqbf
4LcHQ0COTLi3q5g6dhL0RNRakZDQC5IZ2v0cU6PL17jyFeY7wVXRMFy9BxZZqgqCGvHMNF1HI0Bd
cKGuqACf3i9lTUnqP0AliFLJCAb0Q/gItBSFgfaqnQ6qgbltPrVjLF7Tzlmp+BQRURnxZ5PQQywA
e0/0hzWmVknwFUSVuANeYfe0AKyxvCfT7nYSzpgXWDCyCVttXseNq8QBl7Wi4QFXU1R85mg7dgVV
F2C6Kf3AqhzHcgh2QIJPga3QSA7Im6SHI73OIy5maJ+EEX0TWLkqt6vusZtJRwLKHyqpL5j+ALLW
JKGs4JX5NrgeAJycN2kDonrRLx+DlS4K+qiHfBDhxB4gT68n6ZRiuGyN47NoQpT2e+a5k2qtMbvT
Nf0vMNnZHX2di4cYENNwr3iXb6IOx2U42m+sRlU2Udi/+902OMalbdbGOZ9am9untVRPThEAFLa/
1gmWekbAInfEowJwhpCuRWG8ReP5sN9uLG9hxPTlV29cDVvUqcq8TS/7ZvsJjH1eh6/FX7d48F4I
X8bWYrnKYCRQoK08gWd6xTC3rt+bNZqQBTX58+qolQ2FG5iSdAQjXNEmwVg3sFE6jLyYBaBlXJ+y
cx2UI3nvBjFIkoO/3wRA3UovRijKWlzxEowpb8fgUbkdTpSEV+UyPb2TiD86uwSqxJxXh7DxAHpD
IG0pccjopsp0PP1qDICyVraT1rMDziGGFaJZhOijyTeTj9kGZrldHexaU06N92w12qOXyvrVi8By
eeqfygAw0nUkjtO64Nze3ac9AblBbn4UznYUd1YvZYfnCJ1ajFE7CRfkj/5pHrkobA9T6fMGZ8iB
eld4un6b/0Jkvi1jMDRyzRnXLfZ/Dgvvd15aqWd4cUBmQdyMaqzU/4OfD9vWapi7fzvTbMBZSSyb
U9c15HmCuJazCWxYlgBlqEZV8M/RGYHijaZ5PZWzkVu9wctXe1aj/Or7fRDnantRDYDTxQ0p/NC/
mdiykuPdR1G0uxnbqoD46RVLOMnc58QL4apPc4CORwgB/7mQt76v1Q9bdSTQmS+GCrB1uY8yiF+S
b1QsUDIz8BDfIW2T9/nCn/SpFYH5+/1dWIqrTnVxAkx1iWN3wq+krApQ9l1uwcO/awmUj9S+yeiV
BWmD5T5Vjzfh6opFhkQCMKQHpqiyrRCucX2PpYSzjNRBYE0WQ6e1PqFTzkmybKLBazzaw4fbarxh
640bMP6184k9JBLIA1bm/zLMADLorbyU7m9yFZFzrz1cAM1/qSJ0HovoOpvg5bpsylVWnei5/4m4
+++AQM+cie390PRNx9Rpj9KlP17S29FIwdbTpUbXCJKf7jsuMFjrZIac+cFgiNJ4vDkMmR+a2A9p
rDtDrZrpB0OCZLeR4+CFIiFTCyMchBa2yUlbxXC9L+0ixlNKHP1ymuD8z512rmNV8PBrWOCRk+TH
qxAWxiHNDH74/wx0+S8f9ckQBpoN8R/LhI7fgm4w4Vt7x42KTXWsjDucnjsQRs1Q/yUtjLjCZUcX
0xHP418I4nc+YPUi0yvoJFlSB/4SeVPDQcqIzDDNujIrh0khkX6agc3kEexbl17Y0cQ547t6J7UL
NWaDLrvhgVM2QPWLzUQU4EsckfIIbbuyrY/wOW8BlgvJjoiKQ52dYFqip6pvbbosutJ2riH+35+D
PDCj4R/SDSquMEMt6hAdiLqYgYhRsjs7AmPnyE0mjg3iQOL94nTsIVSwHnaThHzKYRsIz3y9TH9z
Jj13T54DTARYqQ536BlBQkuFOwlo1mM9JgdNLXkr2puWNZapLBI9UD0MRNSNo2IBm7x4N7+Ut527
U4YWtgyUI2Z2HMwKlgOm7QY+019OC3MvxKPULdBxhSKZVT44FMMzZzA2O8SNtntKFF73ZMacOm1P
MDH9B4dtVeUfWHct1oMLzHYEQbt5W32Ln8wHeBKtKINrp5JW4Mb97Db4uoj1LT0CRviOeMu8g3rG
gsnnC+B8JLfXMLmqUFht/gTdoL86tGJRLzrQRiIqoX0cNotpaJnJu7zWgvimqNUvdsVgotzfbc42
v1aLW3xAYuf9Efg6OyLb2uOYsR4/4jf+8l+RmSYn8y9BI3HIlY9B4Po+ja4R1zWP9K1bPzeIad/v
Zac02kwu5ydHOnj/hZg+WpshHzHhhLVD9pvLdX53nH+BUxB2FYcG/ImCfOoQ7p3T12k44XjsmChm
n56ItNmZTQn3oimYB4WPueE88c+AOGRUh5d4A6K/uudw+AqC4rIMNKcDK5v+rB7Eh6QcBWU34NC9
3XzGCgsHtYsniPBW80somPT3auFm/Wvf/BXc0II180SI2UWsiHtZyPMlXUW703Aok8ypPhZs+44E
dr7qmN1ZNmFlN/tszhNSmWNLUXD4Td8VDDnpM+/jKMfPJoq01R81Gf1DynS17yei7sbXx/bqZdqN
yWQ8gYhrDkJb8JVysFNax3iMWsBDRXIGgEsbT8Lc2EZVMaKafZUqzgWIcWoMpvQwB7sEoNvAJEmz
Juw0hJIjuHpSj7gt4doVvMsTXRly3geN3SVBkjGFsiiq1PUVvvDOUtGeEADrgG0oqJ5fsJNa/CiN
NkKCvpb6GpdFMYruJDSW+8tHezp4ll4yknLi0qnloYMjNNSpCpBu5DsxZoMOTKPIjMYU2aOdiqqi
M0ppZ1KbQN0Us6sb+tLhnV2Bu6LmaA1UfOTEDKbxV1KZnncWiUuKsw/1+CJgCiK9rHfYXptOPj3Z
Y/cy4jP10M4P3NhbkaIbG2Rpwyx7X4qLULcjNs8uTiTlNalae+d+zO9ftekUWyOzvQpXKALcwoj7
y11youw17R+fk7seRzSIrj2nwNJBTJ6Oq+A6aq2kuTJvgeTloMmhaTNalYM9nfewfKQA4uWcQX2C
2pk+bGmfIq8onjgt9tBR9IcHyaKaAPG9S5G0mbm5Qy9IQpje/NK+msPqdyhtxWdR+TjpgcxvP/os
ueqEehrM+gEAOXM1q8IFXy6sk+qr5Mw8PG/C7tBVK3q7UeScucrYdi8sxkvEg2veIP86Y2k6QFmd
ta/ROfK99HumHSDyCspqaFWWURn/v6PvthAzhB/osJMLeCgtgJ1c8XcRNlqUprltkxOARK/V9OkI
DFdqYAx1m0Hoyj/eMwNbaXnb652O2kHefKWdrqk0HSUslJa69dhjSpsFHyewzQjMlT+2ctZA1Rku
VZE29hX8PA1nma10FBYG3XxaZV0hOgqP+9VwnvEvhYQeRyVz1F3WMbBa5Smiw1yjaas65gLx1aTN
tGxS89XRaJyH3G3+F7Jf3CvFnw/eIs77E+mrRM7is4uaORw5YRPS9JoMUE6oY8FlceSlq3vMmw+6
nuz6rKYmGxWBkTLN4OPZOmHvR704vbK1te6s8apTQWFdCub9tHxLX0pApi7ReLuCBT+cXpRsuNM5
nuAqe9b2+kvF9gjKAkemE2D91txCx+gmRMxuok/itZZ87UNnjGhAJK6rJmm2VrAs0QbePbNrABod
PpXsn6wqc97VwLmvvn4dv4bMkC5+R9SdjBRdj1p6hN/2o1IS1AL+yLkpWYz+a0UEkRDts5HeIGEj
LASPS1OT/EH10MyDjX31mK0ht8s9ZpdkuNLtC9lpmDNejyDMMIZNXW7hnTibjy4+Ro1TEMplqzej
IagvrTbVYSNf0ztygWZ6R1y7I+NC/67W/tbpn6Y4pddne63wf7rvyavg1+Num1bZaUidzjgSDQEf
UKABPJHCE1z0HyfSuABJUa0osd//sOaIP/XsSGu8E10V984cCmf28393vcDwzDFH1Z1XwkmeALb/
bep12uCYpHm64MKA1Du5RoFelHjV3jBsqeMBzgWLnCRmMs25iwbSSLBpvL1xdWGdiNhn4bUVae//
KvH6L9W02CTKGQm9kvaz49/cNquFH0KaDXLUR7PwU6TTI55a/jy+TIk5q2OIwnshFAXh6YujLL+v
ypBVXMlBHzJ4v/8jYG6FDFajsR+NK4rZkDms5NXGegs1fm5ISEGGpiFUyOrVipgjl2VRSA1utwM4
mWhsy9SYfjv/EzlG6g55gN7f2NLq60cUxSjiFLU4Q3BjA6hA2o6rkFvtUnd44f01ysP8iRm8AhlL
PYlpiL9+5rgKteHZM+DIajy5dPrweEzdDwMyuwSJAGkWs6xQcw8sIJygWF/fVsIpG3r+ezEMNeJU
N8wkMhQfzvo1KYuLbnPnlI9WdHCjoBMITqp6fUe15BZ/IDScWb0jOKIhq1NZLY2CTDPKmVuLEyBs
vfINNn0d1xiMjcAsq7Dee+f1st+bpjBZqTFgyPA4YNz3e+HCjtEHWyHMz7XDn0W3ggZe+JP9eFFk
saCOalHKYjZB3cOQoaGxlq34SuEwv++CjeO+gax6zhJ7HyDUwaiigEOP/hDwpKlPCYO7ZuuzqKbF
KX8JC2rARAW80jg9SuWS8dHsvQthpwMQYQjYnSgXfRRIKHG58j/Cmlj8tfUcrrV13P9PYsNp5M35
56PItKGb4pqHnyIGu/igFOKx3qOjU8MIiLC3EYnZ/xnGtXsGBrJcTkGNV/VKnXw7aHGPtGnYaj72
ch2u4LJ4eFpJMat1wY5/ioaPHH8I7GC6v+tnsbG84ELAUCwjfHlJsRxobkSM08d4Sqi+u52Jn5mM
cK5wLg3tz5xASQ8jMb48lQwcrSleTV4Z6kBXqoBsv1ccqt2fKSsUGF1gLizCwu3AT00H1mXP5jg2
9q2LDdDQoSGhdRLf1W523Oe14PFk+sVZYiFxVJyFcG1snSXTJZUeNl5Uz1WlRdJ9uzDGxODMssEC
luHpN5JWeEVQPs6NBzPMh0MCNd2hN2nL9XTmg4GVBhNA5A6hgDi6GjnTq9OYOdU6JsgXZjinA0zm
SlqLKnjV71KlrT+WQZ/PfbokCmd5KRCoV8wqTT3yEExH9UKn1B0S6A0xRzbEy+5IDd0RYRJDkaHF
jL96V5ItvYwFdO3X3AInCnwkINroklM9wuDhHSAYlnUSRRnJ/oAsvS1uPM+Wknz0hoHz4PiL25Q+
q0trvGksVTiuLsfiLV+xtqJQfzTYj+QL+Cg78RLiTO/lKIRqU6Z1JLRoXGlI0zv6HKyJbzROmv8B
Dsn04D/rGj2YlbZBa2yw08youjYK5PKR8FcZ/oHcF2rzL6zBvTkEW9oZMPhXzCxF9DWXuNWKD0CE
EBUC6Z6osO7swoMuowek1e8VXT+hpsbA2gwdm546tvmHm1jMUi/pYEPPd/Ipk7fqXO9rZGV5QqTf
BrHQqUv8luYce8KGBSqN9DrmqJgIaA8obJlcgJET38BSgTmJks3X9mQMnqWSdUuvDse1dHeQ5Rwn
Abxm1b7kFaznabdd4AELITqQLgoiFKyNJ+EIvJ8sm2eb2S3XYfAHwitWWYTfWiAznrTErLVoe1wJ
zgA1AC3+/SyP6x5fqBkKpXcmHM7KBEx8ijFLzlNmZyfGgZoPwze+VAFZ71+Sdh33CmzAxHzLhgwG
MKBUOXSVNPEsymJbh96G8QKvktb7mpCjzdleZfvqW4eKp50xucKbd0nveO6DxI464MMHOTWAMMde
QlCYKnW7sfsEBqrzwKVHwthw9z/5wrFHqFMuDRP55E3TOZKQUfSGS4igkjWktRClhgk3DgiNQ3eS
u4FFlE3HGG26CzRVA9Psw5ZkKacJw9LYJbslj2lcTu1AYOGLdGwHs0wiKDCukUYK6Fj7OnKA8jPn
sW3qDGW7Psi1jvsvpu5lrim2OKlb1h558MHiS4xMDlGU6O2Ga07FvrGo+hP/S4kvcwdCNiFawyop
jvqlSwg2cCViZqMhJt/qMzBphMu5S6KBKrnv8nP2fWVpqzzxrkEyL7x2jP2sriKbbKC1/rQgzbZX
ByKIOyIB3qDKM59zZUAZk+W4hG3PrI0fjlLLnJPgMpXTXo1eQebmPmJoJ/aHSoGQ37AUMveNnc05
GTpo3gNokTKGuQFouHszDL2Bk2No2Mn9XtxQioY0F8CXLwLBbE+yC8KRcCklDsfKJnfZkKqrOqG7
QcSFKMvWYj3uIaCo0H+VSD4KFOz9yMmRn6xs/f6CYCjU07xuaZfyBwpvHeew0l47AmG1WY+AfMlI
xFVzRyrj9EWoh0DQoKyDP1DUf1af8RWPUe40indlJsb4kXRN0o7NevOeO5GcXAV6lo5RsYNsO7hy
e64Oggxa3aqX+y/ui7NdSsFV7uxI5hqnFrcp/7+PVy9buMV2VqHbSeMVfcqrmJVe+dFyz1NuFn8n
a4I67c9UB0pWJh3Y1NpSTDXDX/ASV1c3Rdif1w17GfYfudQ22yW3f7+IORw1Okj4a4uJF6XmLrmx
+TOKoeQInVZJhSUZrfROyJADz+BsWjQlJEVnda4fIVTx7DSxdYPpZa0YRloUA1RrRloK27ruNLgd
fAKgW4kZYM9Al3D0/KnH3QmE4fQ8VorECgjPAKqByR19vZ8IFsCVMwUer8fQTslDTEH3PD57wG+J
3g8cplDFtFxAKSiyJKk0/Ym/+wUx2zdRoyS4gi48uygm3PbYL4QWobx0yde4F1aKBGJCoc8PGMh/
PtaUisNGuOnKyxHlGyrLg5jn85cAWJz5P8tats/D3eLUGHmRi196VCGaIOzk6FwgvwHKEsf+cPPn
UbiDPWLjrwCmRPhaThboJUrnYxyco5NPSxdlYfq/Sf1CB73qwIAtuWUaGK/qQFGc8AJEDelFnnm9
XIDLihJu+KwicnExtHo+0limHQLmEbLZh/NhlqUFHADK29CIB+PFtktSbiyPMJz3Aq5ECWeOJ9x6
i4dcIRM+gibmi7GZCWORbyjrK0FkiVVMuJo2c5LLIdkYdR0Q4FQdFM19gbGnRFPAen/2UwW4e2Hq
hCKdiKOX/4oB3Bm9GZcUGjqC/X2PKCb7WjxBkflTpfGO3NquGUxeCFrmas2Od0TYv+4wEJC0dJLC
HZ1bAmZ/qc4SnYo+UJuyB2R+W6wrrGisfh4xcW4tkrVp0bbUzV25SYGrYDgNF5MTCoUpKvGHdF1J
ny2usyEuxREz2yGYzG7Xxce1ZrFginrbPs7AnktoBa3VAddN6JVVDsfsxcHvvgT7gG39CcrfCnwn
JYw4eMO5B2uLqLwOa0vN+8qfTGa8oAw+1UW2sH6UGTDhPTFhrnQwAeJH1sGuLIrbAflWUKE4recs
5zEwOWjsc11PH5ngaaxVHkRh/9hL+ciOE69dYjxUXQdMVCMMOqAP6/7XYJrNLgU74K9gFxjWw2mv
Gb3fYz7IumTCtfYkqSsGHDRnwz++OTTi6G7PUvmYzVUbTqXiL6ewkkA4nuMThuok9LtkfjRy+WXw
X50w4a0/7KEWsjlSjfgrDo3mLYNcExOaXb10U+cH6LAi+6F0BbjoBhiWAWNYkSnpPP/uEfM09FJK
yFioA4WKaNftZV9FwzG8KAVwNeL3TNH5OKEuUKOcGNBCE2Tgm6CMPJZz8VyMihD35MGHdf8JJH9f
K2SSaNFzfvFqS0A4FzqbY8BImDibvaU7ljDHfvXryMmiaF67ya6Epz3tTdioVT1iRCcGJTH+53g1
DdRyD8CQHt+fgSVNfOos859Mm3z+RPyuGAhcg743MVXs/BdsiAMHQbPQmGz9ZqlX55s25vwANefX
OXHPitVl6mG0ZSy6vbTMBwJClxYyhHAwkt5kT5urNkqWPfRICVJhppkw3ULB3dWDyn4NRz31qi6k
oU8ugTLvSX3mig/H+F8ddImPlYvWohOq2/uhSyTtUTM2QPVdIgWklKyyajqrlz65WOrYqqDXyskF
SwArdTmeiAY51AKfbWFKHy9Z0+MPO7bGBH1/IGOGiFjZHSKDyjypUilrVIS97M1hHgMcvUQiv8mH
4AR8STn3USI3G6d0hkSG35NUWFetC/q8Zs5Y86IIYoBgDWNyX+Ko+9gwIRolHPDbVbIjXQSXFhfT
BHHzpEAbD/qOMPZ1F10gvblg/jJ7Vgxlsnr3i96HfF91Ke1vkNJADXN5+/7e8ScLGKVHv8OimtHl
LQ1BkojXXQ1Vb97o/P35UFUPa+tDfizIzVDQbMpYQIqvBOhBQ1ZYg0tYRaHTQCPymYYcOh7f8ngf
fW9baqbNci5Zv5Lw+0x3tg4ZRhf8MjvtvydJ6qXZhT4chkj6xm/MWx/691ATItXzx0A7wMen3FbY
NE2C7nHNJ8ee5GSeyR24i3t/wjVEzwlciz1e9XLN1ht3YGyJtUoGu0vmE3A3swxv64XpibB/i4j4
pMTks+UDFqVX9rLeJ7JBP2i92o4Y8gZZ8N8vBd5ennfL2kPFccYEQLplOf+QW2wwIIqdWVJ77Mg0
HLbXDSjNx5wXCaFwowcssQ8M5ag7X1Maxlw8GlHxCwkmZGZpJzMUhDpB/Z4WwNazlrcSI8H47EK0
qEMGcyNB/XNWIDvZF+CHDgEJZEsCCqmhUedySIv+70nMuDmHx0Cj55dz3aauy1Q1QJDX9TruCnTI
+0cErWGxRj2UafTaZW1Vf+JBe5XzXXQ7goZO+EEiXBZEzK9CgnAMXys15hWPUoKuaMsWFt+xWOLD
6Xl3bqu2g/e5h3PX5FOPyQdbf9Byfjq6JmnqFEsbmFMhTDzKPBFGPe0aACbSfLUR6bRO3jByd2qf
wDwubNplP+hRFof0P4/AT7B0ely3PWul63eTMwgCJs1LIxsmCQZOtfp+lPYUgxUsPH8q9KCPaKgA
Sxl+202NN5+on9P7V8seX0xWlq00jzGeZ6kCyapb/wLqJ+HYmUt/i8n4FDvR3NJ/PoiR+F/w/2Rs
mn+RCS+L1NlYzLGi0hXG8p26cZpFjljqFVIso/VeOK/iw3E1zIkQObnrWhnRyEZwCycaUXFVNKFj
b6dLtvSG8OxZMpKyNBkoyn8utD+dvIXIhVGCJBAZH3d/zqto/BtNKebwPos5sr9xjqy/FDJHm9En
UaKoWP+StFLHVCPnET3QOQ3L7/c0N2he83ZZIV5FU0pDUsp/N90uTY8f8eAj2t1sTWSYVRQIfBe/
z56UFg8XVm7rb1ShAV0+rb6qLJ1XpKbjKccQUEFl73vf/y+ButFD/jbLsADrkTuqZVYjpaIarJSK
iKBCARPsDm9Iw6HUqGQMhHllU9HKRJ9WkSQJ64LwPq+9q4u3WgHFFGCkOh9+G0Xr8RgY77ry+fJg
ZFkFVmadx+RVs2LRNj8jTFxoyg/OGTdQVSmKn/xJqGuECK1ukCwqv7GtESWVwpOULPI397f9BSaa
tWaklJ8R6/ogQQgtCE71CD5E1ZWGlFJaql7k5QxZYSocLc9QeYmw1Agy6PsHVxemYG5fcqcG09Qt
8c6IHLO4iMZ+o6UtlAPGR9s5lPrhqSnqcK8AEf0kE50FvP6Nl/V6pLbormaMESTMb+Fv8W0YBSqD
H3fKntI6GcNB2NUfCs1TeuhXn69SGowGTbTt9AdwmUOCVlszMAmtG6cDno6WzRY5381ZImJlJ+Tn
8wJV013yLkQdlyTtxIul5GABd7NpEVa6Mf81KW2V4DNoiP3i5KuUjuC6YcmWKpS6cmvm0pkheNyc
jNNYJ0RGPXJLeoMUGEDJe2wkZUF+f/lK48WKucleAK5DDJDG5BZ1OActEbfKzNtCv5CVW7pocqNp
eiHQVFvk9n+Al9Mh5AVQzHR6bVqqMJJJU4uw4EyqPAAfOE5aHUfGV35a4XJMAiy4AYHOnaDYG/c4
00O6D6XjFTTWJ/9TySdGITGnkobgQnvO4lZFKX12ihAhy1NMOWnOcn/3wbXdEuv8dfn2sbsPhyI7
iWufvPvn7Q2EE39nJtF7K7FUo5qqma51kWUM2g0uSx7/U6hHVu+ixbotNGUY2w18zbZEUr6/e/2f
gm7kvE5sOf3o9cJfB88jCpPETnZwryFDuUtncJyKa2PTGTFCIF1JIHWSQ/haG4d+7b9wTwsW1jVt
80oy7GOuecqfnLML6uaj+nkvnJ0CwRfTtMr9ZLQU6K8mv0PPxR/kDmvf3c7E/CLwxb+WOQtCZrFT
rtyaSrb5jFPuRkDxpY+fXOvePXxwW8k8vE5dFS1LfIsNLrZ6HbRb7ijcSgd6QxayVyuJebOmDqSu
QkWyslBqfSf/go9XloK+Mx2PkXAbWo2bGnpXdAv1d6v3mvZreRRvdjqJdf4Qbk8tNRf+0UzdNr4/
yfQXVIAvrzVaOTAARB0P4P3qWpkCI5ydGsfLxWQjBDrFOBkcxe6RKoLrprGeFKMhgsznU7TE4eDQ
UcGr40kiebMY2aoF5EqQ/k5Rsb3rKM9/iQRS4nydtoR0kXcYklTNtozxQc0dtV0k4GsSlcYqXPhg
c08wy0XQ3EVAo3eLb7wgO59pPM1bLWBUjREGUCHKhj+T/B5+61WHGZRjrSxSaVazX2Azm6YMEr3k
6/Dsgg+t0c/+iFBTFD5+a3VR+rkObz+Tuq8iZ6aILYr6f+uiulvGbqKSLiIN6nDd1RqbqZtk0lZV
68E2nseKRdTlpKKYftCc1FqH7D5nLxo6ghc3tvmoI4UOhTwRzbkm6Z2xhXcH22lnwhTXhdlsMuny
ftkFMk4T2JMH0Kw2kfd3AApvtODMyzhdBs13kLjp6TZAYcDUrLUfXlRuxGFwYSGdZ9ppUakt/hds
BZ6zChvNexsE4+Av6kCmdJxbiWAF/CvMBlYf8camozvHY8lc94JL6GkKtLdKpa4VtLIUWbX67Lxr
bST3231x5M3xrhQVbWzh77MuFxubm4X/VL7Ptj7//t96nMwZkq3qxzcofp7rukDzU5+xqUQ8QaSa
N/YIi7YpcQZ/x40129MN+p6KWR2C4QFVHpIoos0mmVngx+woqA3XJGjzyyOqSDtscrKG7zMgoxfb
UGf/Xx/kVNg+NEZAKLteHSf9ywxnjrf0r/Xl2i0KhvEne0Vy9vQHUirlV/OCEM4rlOKHNQ/1TtRw
iuLV/QrAtdmArqb18C92uG3fIgmyCCYx9uWbIP225K9MFBu2YadVwA5VIYfLlShFd43eLTDh/XQJ
cMcp1mKihs2yGfVAJ9b98T8/eX8RxOe3uZYr1a970SZB8Cc5GBjBggtZW4FXf6RmhXiPx/AW8wpt
4kViC2nfxyYGHEegsXhU0BGZqTlEJh4Yep91MU6/LKGkykWwLfiSbBI1s05rxujDVIvk5cfbCXo9
TCZ4jO7c9Ti0TWDBK9IcU/2EMbTFbO+mrG/1zY0SmnCNqxFRz13DQ8jznwR6V0OEzL+UY/8r0r/b
lu1XUA+HV2YDFnteS8hX6hgBxeezYPG+0A8nIDbktDWVnetUbWnahfWaqBV4pMlqlT/2eLziDwm7
fkRTjScfvXPWPSX20+UnWg7ftbz3XnjXqe0HtInPxNKXbh0bodk4RvORMFGSTerO0MHNG5vz4FuK
9DUidlG/IgD9K7jSbsvj9u/hzvwPue82cqPig2P9Tvn/dcZFHpelgscIxE+5TucNIcgGVu5ip6m8
tEcssx5TJYVs6QjC0ak+EetD0wijSlpcISPmbrN7hQCE05cu9D3ceknSZbdmzHRPyhPF1+dRP9fa
uGrbJVLOUtNl8bsxMcseaLQF+y3WvOfCZUiEmlYbEKnZGAdqwk9SDv9ZZLX/qIy096aS8j2ff7Gf
lj27Co88yWlO81MJBrMHNkKO1e0K5F3Ypigm69KrZ6YSknBoLPYAkPWffMfYq5Ya82CXLxYx4RhW
7nyQlwoM3ICwSNz+WfRTErse6b3O4Ui2qHXyaLvYqmhQ4syzMamlAiBzTxcFWvimdOxbPYlyBS8w
KzudXiykYY5jWhSoce1EQik3H7YX8uPnWTKcVXdXS/VEO9QKV8oOeQkOBXcTQYk8VZm/jpW+fxDF
QSbgC04eok4vPyuq0OaLOknn2S/x81g33BvQL2UVqbOW0RugKVIc8CaIkzaBC7P61hNonuL2/Mri
gz3tLRwIjbmqDhLZxCwSqGi9PeneDFVs3PeTyxGN8CwFaq+QOnZOMQr6dxo9gklCHUrl1h/i2cv5
m9SYXG2c/5I9m1wMdXzClfrwleagIxMIug/NJH2VmOnbMtAz6dhAgFIbdda4m+dmsAwxjio0oGP5
XsUPGFh+y8pjR7VNxj+XvL9R1f3AwqvN53N8dxf0UTxhvFNyyk514F2sVGWC/wmo/2KUGvFY+FCE
XL9tGGe0mnYuHNUYCAqXGpeh0/oJIuZ7O5a0aku5opUvBhOo0H+7ChaHpYif3vJcT066zayguTg0
Ks2SmIUiUygctpF4TGa3cYcKSusEC/uA1iO5Ps5QKg6ru1jcU8xX3shjVoCaKJVN+H+EJHt4U+uj
asv59DhhJl/+at4OIZWMfjRjeqVloeJYdLX/v5bFIcsC7oIyS1eYBjwTC4JkaT2wxUCoy/hI+FYx
wHJoEBuXDklT25nq4FDzdwe/yPfHECXlj6TOugbxds8n0TIHhDhgegZeIMhfJXz3QisfRoo4sUqV
OGTTYcywCkrbC0G31zTCJ/pt92HrJu1umvFxNqqMhdPiF28tm3co42TSep4yCst8cVcwEnE2ngCW
Nq1zwfl13JE41pyxgOaf4pi+fChy3zTMYqT+wQeis24WvpIzpILB0NxwXwOeetrodwyNVHSZaeJr
4z6nqxdtobNhMS+3OQg6wPznXuOTXalKStg3IdsUvLMry6E8SBWbc7PJ5LcOJJEiP4fuMk/DQvq+
0RI6MLHRDC21otKdjx+uh/rAosBoOZAVVklrBDbbMd3ZLBQHe7eTwRJm/Y7DTNnGDkN1BeJlQX6/
8p77gPpDt+ADKcLdP9F4JwCC+tW2RUYXecAPVlk8aPCxpg3vFaSUSZayuc3USpRLVvHYjEqQbpx3
dWudU+AY8SQpn0/re/K0G+3GZE0l5eVdFt28klbFstbmQ0r0HEFDeVTOfspYLugBpisLmTedJCc4
Gedfeu6YJBsD0TFR4Zf9BciU11pfL4a1ewuF1eL/6TWxeH4C79l2sdKktS7oiz2mNgSlnz1MAY9b
3G93JeGuKoP2TdqV31V6RIC1O1MsJvgP3tFuYsypXGooS1l+MSszswRWTbsrdn5vLpyf9tqXonw4
i3Hb0Mao37ozaq45MgJ6bMFUgj44yeaVBBfPmOOysqzbkNrbyjqF/LxgS8i3/GHw3Y79xCIsxbw7
C4buPeMTqJzjHkqpaVT4aNp8+SRnBFJkvgp64Oji8toZRJjiXKrbodvgVWZqZ+v7WuExo3p5ZCoG
SQBEDCdE1WLoVabG5eUwXJLIEAVOckrAgAcRkZOJXKE144Vycmej+enCJpcDsvQz7UTASAQUZLEl
N8jfjSdh1z/9d13veCQ1K1Ym6A2R84auge65/hyJju47oV6Q/43pXIt3kkkWtyye/TfpLjX/OOJL
jQWWDlQV5TAcpw26qeqOpe/MxNw6PQkLfhUm1zkZaYtYKH6kFHTMjuhl9Uv0g5v5MaCQ7rIhD/tr
+kCkr2zd0vopVW5lhCQuWqUCvFKwHRAdMHE8jHE+jn5Chk4fNZiBBEV9lKAcbxw6pbkjb2ILv/Q0
t0K87rJ8YfEOy5T8xkwIi8cmJZCedhJDB9xLMj9UKZimC+Rdvk6G58T8+/qP1S/9TtdlWDQ1sEty
sESuuY2YBDTZLiokAt/NUDmXYyx8xskxWOoA5Ut4iOIfEWhjexAFSOCVoapFdCLTydcBj8rGzjEh
c1321CZnxWQOyUoJDAhNfuJ72LSNtf4B+6H9Y49LhOnigcGEjfhye1I+U5N+FAlGZL0AU4DfASPH
Pprh00oxzTs7swUVWP5pdRTxReU2SQ4kt+0GLZdP/epYT9kWoY9hH07V5/VO/tydlOTROBmFXJ22
cvFscQqRlnxxFwcgh0rtutu8i+42VPsC6adRi5fdofqTdiiCV0ZlKzqOI3D4lwAa561T5Dvldxpp
RBF/R4eyDqPcVNTbSQrKm3FC6Bh1yaSfmqh46nBLhQJA3QJnAMztMtNT2kW9SnNkXfJhe4MSAKXQ
vB3ehMc3t2++7dFBUP1RZIS4Gy9T4bhblvOzjCMZ5bJS6n4ZHsxcyGSkSZ1fbKXyQwPiRgDLeZQO
tRNK1jFkoUvQmNAN9r/TVK1RaQzj/TsDIQCow9L83wMcbjum+TQmTz7QTknSXFX7oULuIGx89ztZ
UHNLJ2Oc+E+TUB7jkII8QJ5BRMtPZIF79A4uepqorTXCVA2wCUCeSMgNyjuE/LW17Jsiz6IEUjW+
f0d7j0aJ0BsJtHKOzb1n+/7Mjy3eUPMYhHV9hFq9T+hbei4BgWpUoWoX+QhPhYJz196lq9nIlwoo
yIwIaCFqbSag5nnTUNZW1pNwm4H2kAVG8XXvUVPCpJQFALLbysMxFMLchkFj+GhLWh2yMwqzM8GY
F/1QnyqUuv4IWYogmQnCQhvFi3iMhO6g8FMXnGt7Iyc+NRMAXIN7Wl7KrW/+dopTR47D4hlp2icD
aQuASuIxVtUHEjOLIO2EqdX5YAMQAT5heMi329L1e+8AEMxQICLScPNOPmrbLUtT6zJN83UuXksY
D9Stc8cfoTHSq+cY4/cV4Xjpdse2Dwep3gsoTN6qcuv5HTjnDf7ZJGbJiUzAy79MkGkB2yR+qL9m
GUbzLLxzQRnyZvPaHILMa25420x2oCPHB1wBTb0Jl2oUQv1+eCY/Dp6Q3n8TA5p6PPe7Ko+yM/MT
HgRy9clQoinUGv7p51doh8uX0d1Ty2xSwyBsRDSH8MF+X/2zC+JFiZeK/BfDGeu2T9H4tpdQnIBS
cK2w/2a6yY3zyKZLhJanzi26Br3qINOzivdstSZcjq1Blb4Rqj/Xv4Rti3njyl9daCsiWq7tu094
o/a4V22lvUOj59gU3p5UdZxMTKQzr63AcFZPTL4aQWXzeD3Tc2n6+FLwLMDGWBvmvPJPUW6GIPvX
3X7YOFrzEv72wnVJDXFjeDL3ZtDJ+pj766lzKi21ORxy2YDc6KqQu5DbizMqeOqB4K4ze1NXda2x
cw0BSEHN6Ij0nY03fO8OPD1fhcsYGnTkTyEqqlkxVnSv1cSpaUfJmQfosq5g0pmAwBw0n0d32uHH
gEK91QcPbxh7JscPYltQ3EW9Mzcj3x7gx6XaF30jhM1tiuqA8AKROWhwi7n6KcmdtYEsGqnSokzl
FfoGpdvx6WLgOUFuIrBBOFOfdiI2fgJuwkTWXe7Sf9b80yvakdutkZFF6pIkO1IwJsFy1QaB6M3n
xY3gjaQsT1ISg+MS76K20jhhG7szCWjCaJWkJB1bVFhUZw0wIi1fKpGimcbWF4iLm+NQi0BRZgwN
7GW04ACwIK9a1zkMYDa4Qlid269yspBBh/BoQeHM69fwHDd4v8lpShVt0xfVIXkJJLh2+hVPrWIP
9GNvmtiQ2qIZxFAqlw2FOq7ja8qLzNPvsr4EtxwCjaVjhqQl49m6U7wVGZtmtJcyNyr21VQFdNHK
Lctq3ZIb8t6NWlwc4AbVK+C4kAkAcNKA24D0JsuSAwaYFI120yC6sdp/He41hFWUS0U4Xm0LGO94
K5KBsmNBzDZs13L3bbkBxY2g9KDoiygwAHtQJR7ZIqn9q0mK68ydQlk9tZzkO7npoXTHutGQs7sP
Kru1a2YII+x3HBuxJqjmg1ZtbkthaMOWbumwJ55KOwXJgQVeS6PSlrolQ0Pj0QPnwohKXze7n+zi
9L5my/ouHpCfFJun2svvne+2p2ZQeW5c9N/H7I9DJsj+72Z/DqlhAU3eF0vDUevEG/G8m6W7iA6H
7aKOAlwWGLAsa3bXeBGccUTqX1mmuCDt3J5nGVExy+MLuZ+vlQuztJprMwo6tulUz1TRZH33Nu2P
KYn8nmcMW1rsIFhMhk8mI2gmP5fvEM7+YYCsyvE4fOCpJKzdne4FL+IljQuOogJZ6QHLU/CE4MQs
e5eryqJuxamMw/p8FarRR6MB5z9cAG0LGSGP3rY1Dw7zLddlXmXAwiPrvumH8DDiCFl7LUYGEvPh
oiFVzP452kpfuBIeyygJo8OJASmSCdIdPrWCPTk8xg2E2YfA8PBVx4l/WU5lVOviPSWjVRzuoI0v
P+B/wznd60GJRnhC5llT1E8gIHs4MbxPXs5RzRaqdqrOIuZH8/iPEuBsPpqQusa6T/+SAgT4j3CX
IPfRqei987xYGrS3IcQynNDf9OZ4s0Cho3FogO2anLNH2U3NgdRh2AOwrOkLEwnyrxrfpN9BbNnU
UOGfYCLkkRxs+FgySGimJvOOEKMI+2N0j9oz1Da0yQGK4uPay6rIbDXxlmNbNRmNBY5i5Z/h+8ER
eIcwO6n1VlBe/sNfDbxRoRW5U3eQzsnX/Fu7Q4Zkve7g8Qcj+PG8Vd7k2opZgH5uHOp1fy8yTnQF
s6RSihaz68BCXbCWqmB3oNdoSie+VUtxzBSTTjmDa+oCrJPnx4rrKRqlPKUUC0e6l8tsE+yQ8BYO
XLmCXHeaCIH8QQBGHGsA2/BHT2dxEgwYJDT0YOONvF6nHUkBDD/CBu/uhdvKckisJbpmn0z++Q9q
MMEdfBcEk7G7NfChKiwJAKusiFvkXuxS9Y2w0DT19Y2cxL3GFQx+/cCG/Fp4b2a3v8d8/BjQdcUP
8dwtFp6UR3F9JULq517yRNb6ssyCDoCxqplhbxdpo6Qwh12NPcmKlbHfGAT2v2xEa4cBaWWSOitG
Lh/SJfOgUtNzwMHyl2LKRRuPY/BJQhcbDUkINq7g9wA+Q7jYXoPh9oXsYeNZJw00pNfCSmuQqeAn
b3+98qTSyNt8TOEmyMCJOBVgNDvbG1867uvpWwCnp/VD+rrXjsUCDLEIfX/+J6a4iQ+5H9GSp+2A
HQmP4IOFJeZdWTSvQIUQvn1osN4sdrD+orfaVzHwS6vBeHadiJir9VdezmkuD/vYMdnHKiCz2sB5
ZyMh2mwpF5aKfSBx8BNaK1fmkqMeaXtrwAFH4JsCd2Y9oRUbnrSqtEznFzTTwpjiKFNPIFhP22av
jbYhA/38O98lilojD805EVrfSfb/vBhJ9LrA6LWQ6qCVWqd4U4oUaWU7aEaSZbXqLUNdu2hVIMiz
oCOXpIXlKmNdKEZe2SzsEh9ONkvHxavqTGT+YUb13LxzlAQNykLISlbiGVEqnFqh52OVrv3H2/yN
ANp9dtw2oPX7cWobLt7lBEk8Eq1Ip/VpLVLEZgQcAPR9Btt7ZNAyBFfopMosbX5S2F6Tj2wYQ8m8
NAUFPCFD+rpL6F7QHPm4viIbhZHQZDfbc6oSWFYh7ddPFLKfdQuWThaRZOEl6satKlW8oUURQ4in
BGYtTiKwizHNDt2dBVobczn9Xxx/8QZULtbJQH9VO7ubdX8YvkPI34kwz79Tlnc/hvzwTTduOwmX
7N/9US5OP/JhZN/JQbhbH/QB5IhhSvlqU9CoyklmKAjr6PHuzs/vMEdslUXyCzik5Pku5qyh+XTX
kOOArKnG7QC8lvlQQNqq5kWVCR7/nkGaM+u8B3WVgCj56Inp5fAwDKDFNJFlL6LQ3ojQQ9VcM8IW
iCp50ZsgGSwis4kxtu/+htHWyKVFfAYr8QM9pfemPsksK3dIlszbmhMb/2EeFzMqWn/SGuSpBtBu
65RFKzpk2I/qxCWXQKb4p09yRUID4G3BrEH0nhXcIAQihffZgjlS6wuvgMp6XrDqjcM99txUVZLe
SOlJC90aRliD1N5tnxyLxeg3B5y3mHcTDi7tqxMlcD5z9gG73F3tnci2ru8ybJJmmlPuvC8cO6t9
7YUc6Z2UZH1/XXFKKg5Jf/pmu8k/WGzvmDHcXcLjBj4S3EipPTyJPBuYgE8GECL0kClXiUZ0J525
/04H1V2xBMuiABRiLxM9fzUHJVUZFlD/MmOLPr3j57Es/9n7QEZxyq5bJofQMFdGD+F/WEXrqfaP
tJPuF9wcGNIEvCskjOy866p5wNTPuqFJrmelFxFzzB+4KCO7jm3B7AFyoQyb3Bx/uLGP3megJWt4
fVX+4tQvzEcQzzmBMkvMPz0AZhiVuGgg8r1wp0mX8eqUACFDrtPAmQfPEwwX9E3z0yy+cMT2d35e
n0ffBcIy9Slo2erGLIL7RWv3wh+waDmAC75Hdl4mfLlJo26qf7T6guxS/nJL8JxP0E6hDFRxJXbA
MQCbnsz9WQMJvinAD6ggH9JkSClB4DnknKoXZJmPJe/ZSdP8laxPfEfYJCuVs6y9TtlbeBpUA/sD
nGLGLKEVllELmf2PsZDzhBaSuvYByNrig7cmi3P4I3VjFU85ytnKFkeyjl1K3+VAEDe9XmEN0c+/
02uzH0MOXhkNC1Jy1vdf+n+YbktDmClkbnF5LzNqIFQQYlfH+ZHlYUoTN3w1oJVhXvGdC7ilNFkF
DYIUEP+CzHalozf7gMHY7tEyyHMNsp2XWGkngdu36tjDVvFXnvnkWISU4XPbU6J//r2x7kLG4YJP
PWyVeHYcikEeu//zQ7fFtinbP3AMgmvHG15DXmUtgb1qc6kNOB102qTAJShYWkom3XixuPz1IZ4B
NjtprDVmoWb1+l64PtDp4+QQkyYks7isQVdpQsieMnW0bxIluryN5KBr8GnPXytpigxcQCDempyK
nS/EJGS2rCWGjfnCqf89N3Y/9/JOpPGVCZmkXk/9BlVeuPSteQzfvsrEr+Oh9k57ZznMU2KNEdTM
m0Q0ZLuYFFq9xTLHv67QHOsaKHAP2q8RIx/W+wFivHZNe09xgz7q6AMwnmj88Pjwt4ILv54jFMLm
Pk0liC3NJ/AAIdX2Kex+x/ndejRGs30FXYyQmnCxXNCmWZqy30WY7nMrCcOiOCG1uj0LZjIax5fb
MYpfa3CJ+Q1oYLsXFw5JTHSiC44FA+lFpDe0MKk3KXvRQNyBcDNjPh3k8ZaaRBaJnH2fFYNePuoD
tyYdiXB8/WtSuT1G9At9Yk33JSc8UDOeJUova+F0ifm8uvMIdTU+D5JRIfiUxGSG9JlmdBnQDpmY
+88LvOJ/zowHsBSmbKSdCfvX19AxoZ5er4F7raIXKX8T/0TsUsp25Kl6kbfkAYteJhpmszdGvxZP
4CC1MfAdPcXnk622EvThRQZoCV3vx1kKPfv1JJhREYui6VQm65xHSH1oAQWt0w7/8yRYTXUgjsGh
9qr7NPjDAVyQZA/MTxG5pd2PbuSXxOMFUJSnb5r/vMHn13usVTgR3vHCSrjh8UfPm1WXptAY7Jjn
C15IGijnNs5iv/WS4HHwzFVuhujHVaBl6ZqT3xOWj3vT2eEbLrA1MZipqFXVIX7tM1G4D5fCa4+6
1xcdmW75YO3w6su0mWYtB9nV2XJBA6IeyMJpVN546Mz8deeuR+Nngn9RwpQpXEz5YkitmdTIf72V
RVRfv4xPwaudYv6ixzAh4G4cLS3NB2+rHSOIR6VYCwksL8APle0HA6zx43f+8vsKprLNlePMS0b5
60PmgAka53fZjqGCKnUFBpfMZW/dkzerx45OeFiyctl12gjKKAlJrEBbkpOUU6KcPhsibbQRdJGD
9ryVqkzgUjyPjkrC20GvD9kQJy1bzN1wY3stz7dkL0OxLUayWfL5xTF+VSRAG43E6nT6WJ4Bve4M
QpVu9bvaMlOv9OD6WxSQP3XhTSZXqJfH5tuGfNcj5tZA3YZBA5D978Ym44H6rjQ5QwNlXaFDaVLi
NakpBQcgiepwcR4XRtVCPWsfb3Mx9OMvJqWf7BMZpqzA0YRjFSfuAx4p+kRX5LVhN60fCMbnrRyT
xlORT2XIKBuLA7VIDHQFALrhus6kziD7QsWTu7lnfwEp6eC3JS7jm9dIEser/kiFhGiz5+KppAQi
s6ML1se3tn+nDtwidhYgGXnV/puUR1JVGFr7BGJ3lvvbNPCrAL2MNsOWLiJSk4EpQR+g1GF6WLEc
Sq4hsWSgR8w5csOvvCAPxX3fYblLE5dGfUDu1KIw5J914/UnONBYoMGSWZ8TABHsNRIPxEMh+ICq
4RKBsXwQyKnG7jxJ+mAcSGtwT9Kwz+ey5HWnDdYAQNfl6u7OBn+TvMZTn4XIUYdtMj28/nfHsBfV
9hy91sO7eZUb+xIJ0snXLj/A96JsPzHLEkrFCdvCCNLJUr11oQrRXWsUBZYH8TKxIFm3FuStKh3A
9RA3RKataphZLNck5S4BiVHEsnjNSe508E0SgCfwsgPW+nR2TXUvfdDneR7sBJoX6rqUHSsv0F0k
kBVpXukpHcpTa3uma2P0+UiArM8Sx7GsUmsEBomUXOa/hLgmcGwF75Iojxdlavvq0cwQ6FCGP4Ny
7PnXpaizhMPhR+fgWbxjjwiUrh1a/pz8f9EtViZM8nJzOQyPfVAH5+L0vywXDm+Hx+e6bbv4fUQK
wnq9Ld7DsysE4NiK7XuF6giKDCIlkXvLzXdsCU/fC1FDgT9P6Obulg3JV7A2njvyMiBa5vraUIgX
4PLBSFc3YxrX9qZdFkdh1MKI7oMTqdBq189XEaW4wthHHHf2otynZ+PTCFcCKYAIBg30oTUo6GA9
OPd+QpycVuqqJsHTmOnenYOidFXpI1A1XWriNJ7eZU9NCjixDIZKafAgSTAHAzeY6IihnZQjEyjG
AmrsJxaSS5DaE0vQxCUY+2GoouQLb5f4fEULwetEWihWFWQUT/6oVXQtXV0BK7ygK8RNo+emENza
VDTdWDDl8sspHkGcn3z6CXRhz3hVHKXjGvo4SD1wn+Bds/4lrtCZT4iKnGyGxyr+cT+huog5kPXq
Js7flWjXbNm0wUU83NIU4VFiQROJUgI9WrBt4Zy1FFEMnagjMhUMnfo3Jx/1SPUFQCMpnHc1CaHO
E2qnyeUwx/QV+OHi6rO2kLf0VoxyZt2lNuQqgnexbG2/h+xvlp/1me3+ij40ulkmTvKpBfaqYSan
3QrP8nazKffLucq68Gg/wFxmPIHVe8K5TvZQe2VQnjTFo5d8pdD0YSfPuDoRUZXgcOrXCVC021m9
JVRcZYb5OGulRNLaP1gHAaFru8OrrPwTIXECDOK8vBv6IT0OzRZsJoEPb1SWdgGyalVs6wle7Swf
C9fXYm2HoTfjdiZX3TMYe7zxZRyVQhkFxRjV2/RrAWL7eeTUyKk7jU3uIXGOJJ6VdG8I1eC+F+Tq
+EN8L3kNO5C3E/bFAJhbTqwjQ7QeSVn8EDYrI2sxFyEPEiaMWxbFjy9UT716S5KL9KqS7woV5YCw
G+0W7Lpkj43cVIT2GYD2XUE7UA366ASPdmK94PuvpxxO5HJXxNJoDwcEwWORZMfwe9NpHGrqaQst
k9+tZIMFwMs5Ut4w8xK+6xHe9rxByvgSUazYtbi71dodHr+oK6utsodV4+hz2tFi1qRjSa9Esizf
V85dnj9YzSLxNNAVLd0lCIRHm1u2tbOAifsfeIQcIXGp3MgB/LoOVHI60yt9Afdz8tCWtVZDNZOX
U+s+7ctlWO6yV4u7X1d1+KgW9e1gLh+XGmcNb+0jbITnrAZ5Zhm/8HjxwX86B/hGFMSzNLGYb3x/
8s29+/6g25N8j/OkzTW6OSHY5VkZo5qfIc9a7M2YoWRjUqCpBUScz0Ajv+GG/UzsUITZGZzxRs/S
soGFyUdyhaQeAHIvVxS5ViUP89h8VwKgbR2gYrOoPgl85bPKJg4LWLnk3owtdsfDhFPwrAHqrXvV
dxJ6H9vl9/Ts27cVYsxuAYbCLR3DpqVxtGwf+SXjlIzQgE9vEXdJnNnvTXJpI26CVcTISbgXQpAU
sBjoAGQnuyWt5x/e0jwRdcXi0nahrg6YcApwcUxqbcngsuVcFesWjaSlPtcxHME1SKCelPnLxshX
3Ni7BZ4oOH1kbezLRLfDvsPTVKq4J10x2C/3RwELI5jTTqHN4qkIBfXy8JEvGH9kjaXENOyHiX/C
WsTQsT9n5njvY2UY2giTFtvkaPwnEAoxvxe0aUpWXq0yIx8QrlfxDO5XUJPNDMt2raR9Bt4yrEaD
SlrfX/1od0TXxPnouk9tQHjbMf8d4FRgGF4cXrUoVTQV4iOSCEN8lFPwqPhAhX4vhDMH7XDJF7hs
ANmXLgOtYWgdqWraJY2OvSTtdQh7F+U2ZD5aiTeP29qX6jfbL/faf3OqsQ6YOsYmP7vPDvlEeieW
0Lt2c9yYHPkomczpUS2tlbpoJUOI0MAJwAz3FozOVN+bv08hYVMLR+sth6bUG4HzmJLQfCarAmYM
CWn9GtOVCV/fl2e72Iiyx5ancm/7My7X6eZFxW+YMPmm0eUizPiAuDa8Mucpeq3Tu7eqEHKQXdpm
30ql+39Jrc980MPjwluv0UOCkJSKDm6Dmdp8ENBiF/anfCnlJfevXmMIUszqmMecFG+7HKZNtmym
G4ZpAcWdf0Z74F3h2l3Yp4hcCmKZRtvw2JtEv1fGcsitxE+0ypKYVhpI9fexoNXjVAZjZ3EBLcQ1
rhtTQL/9REbwH50ndgvnq6pgu+2KjwbEwJH7o30F3Nt1kaxGcPv+ASGUqj+zEya0zmZZb3gVTvro
OtIYXGG0K30a1hlKFdUJMjlz017YjZsKyUfOKT7oyX//anZjrDotWJAKmelouleMJR+0AABsEniS
rm+0LRCwutP3/0skKigCIDcbdffSb1LLWuGH8gGDdLhyYfxHapcwmQyOYb5GQv1y9HzNeoK451F5
GbDnIoYs5UNMwCh6M34wg6wKSRgy3BWRnaO2O7Y27/7XWJsOi8ASS96x5+o3GP7ZxJIhI0EaqoOx
BFlUtnxSmv2IFRpLUNylWj66GjY/skTpPzKmBF1KzMAdljuh5drmMsAhEDMM6nAB3wbr/yZW0IyB
b+WxYy19Pt+4FrJw1ozs+7hVL6Ops+WPDx1V4ODvO6ixjbzuK6rArteyCYNIsB4pOWpfk57+gwHa
7DYGodKfcuvXCo/eEVpv/dXBa3lskaglnW2T1ItVI6Z/1DAsXqsl21F7/xjNIfeuZ0yrg92QVc1O
bNXtyPPjLDs10hil0f24IQ+c0+D/NECvqEPRTaCylEd7lgaMyjihc73asEE5TxYVLz3cqY5yObGF
y4X3y/HwW6jzy8N9c7a4nbtc7/BORFLSQl5x+wDS/KcAKw3+y2a9NR0T8uqNcKUgjxQtJarPaKYk
15PcarJvSeK0olmSt2vK/pEFAKDL/Yy7MYiYJ1AxZkxbZFFi1BwVnwl665dG83z2U3tImqLXzeSe
0Xxzu4WNNpq6g8/bEOGnqkRz5pzIx/i4aunn9a2Iz8Qps81rQhO8T1ium+mMtceLnMe1FyqSDgSq
6aEQb+zieK5NURzYt7wSbjWfq3xPk3Rs3Cert/vOSVyzkDiU6/6IbcSc2Sn68n3l52oa8MlZHvwk
buYmRuAiWuwJCih5le5d80lmRo/Gnclzw59GVMo9P6ESQtTPiwSekgzWgtiWxiXKlJArkngmcU99
W5d0yzT63GNFw4QVFcvoZgCWQtxCX8Wa+JY5ovVCDF7THT/GE9tzY6F9uvUwanCSNYqf3OiiWZpv
hZx/5jdBhsES8UbfBGLYdVOfbob2D7ECTFm7YrvzW1lcY5ZWu9p9oJLSgXWS4HEgKsd6W0o3lQhv
wteFWc/OD8ufCIItTDaILscrJgotqW0jTngCZf33T1MUpxXoY85BAZBbOscTmzXcSf1A1DXtlWSQ
cT/VtrveSKN79NRbWFE1mC+MxZYxjxRg7gvVrdjmfKWtKUsQxKVzWEraeI9CvbnZUpKytlXtzRu4
iGD4BaHNSEPqmYJsPgme+1lWXHxD4SqOlnZr78p3kkyX2TmDvTjT5rWnkfXWmTGFWxiLeIAbtTuY
icVHNndOquRKRGFQWRTt43OcEeJvj++PVXDM5wQzQa1iICBOMcUJdkPoSCWyRM8awJBF1R2dCeln
u+4U7haPeFUmxK1nmtDjfkj/HgBp+XA9IEkm9GA6YU3D6Am7QV5nbF3xqeacNWXHr4NEMxWZvGAq
HO55V0EHfSbRljsJISacBV467Ey+CYri64FQGvWz0CCCou/YY9sFm+gSlcqXsO+Qk62IKZLEiuVE
NpvAuFn6gqg1vkbNmYcixgkHUMMsomVUO7QZYe56/Ds395kyrAztsBt1x1CtdzG+CN3lT23Us0nx
IzxKsinBtCRBlUTAeAQm+qLvNBcvzaaV14rCKreXD96YKypu2G7CePObnNEO2DXlCo6BMlqs8uC9
kbcQvQ/BY1YJWcY2qzH0QaxckInSpNQCvKp49qjW33t7AFOd11pbES8Y9NX4JqsksXrZPLD3XWGJ
ex2t/Is0Awm22RKRVr6s23PAvuqOL63wchdvzkBNEpkQLOEj1o1WT447cZiDKsUuh1Rcbe4t9F8B
xLSJOlOIkZVKmfi53pJxMRXH8DSlrHMNv0DQg4eKDqoELIoiCCptkdkxuR0QQReUuxqUG5oeqVI8
/Ra+Hnapc3oaH0YdIy++S6N0a9g7zwGRwlGLR9UJgI++AZUQhPm+Ohz0sQpAw1vJXJTDLITBx+TG
mizQ9aWy6TzLNjAMg0TcHummj6ZP64w/0mOXBsR2PjBXM/cHHIOvhX7yHBm+WchqM1pN6BgtIcSl
wGVEdmjiIAdRsB/hQn/feIO8J2lcHiiD2BmFikQkALln07GBrNB5KaABqzzS3l/s8GBFJ7DH7N0D
uFvRVC/RpbWd6KDRekF9PaVRtWdYgPJJ/C6F/c73WiIdOptKOy91m3DNDXTuHpmvQWc5lPhiw1Bq
alz7Iv7xtaDVH1G31CDWpI+A8CHDyYrMFbEql8E0FU5g9mltnIkYYAjRdb9d06CoqY6mby49RXL+
XjnDT68VWdDVdPrU8N6hj+pAqk96sndyVDpihrCGg0MecO+rzprF1HJU0kiZP6WjEUzTbFH3x86K
Y+JAyFLw+MiysG4QS1p73pyZcbo7VO9dVAJ7TxgMmKkTqBYvgNmlliRE+surLeXwAFThUkEcfo/f
Dk8rFU7V8zBwNfyIhnEY/jK8VnbSKbr54Ccq8h/ktz7mPkp3JrApzWPbRG2FxlKR189l3cHSLst4
B4oIrvh29C1MPtemfhAO2bvuqqBd6GVssauyNa14wusb8ECbqL5G/hjsF7MRJvER8ED2AA1yxoXx
CKXX1xn+o4esQzxbKycXm8QhRfYFrgdhR9HdFR+E14kEag0GfKdegNP116BbvqXbRE6FkLJMW4fk
bFDfyzBB6o9w7tCmAhyjortaMBNrZb2EhnrFRIBTvWq1UObqKQm05Xb0y6YS0GSEzH6lQbHBjuje
zh8utjdi8+/bg/Cc+CG/k5Gpf9X4pLqt82fmasCWZeN4i03ehgjpReg4w7CEF7p2IzM7CzJZVRgZ
MbpgXxHHNkkcy5fUE30M2cWzc68RJaM7hmzjoXrFS2Cs/bQi1RWucVZoC6TiyjVcovurkGf3g4lF
q3TOzFN9q3nRhgp7aDsjVkfMxF0xoQBhwKLkyCgpYXhwmystGPkqpg9vMvfXpuQTFILzLhmDmmip
VL1CuDxNDzyzfjKUitc0bxekP0hdrRFiMI4oF3otBfsIzlKUTZLxyt9V9W5m4g7jLHtLeE0BWqeW
8YMWOwN9kKT+3Rw95HYFSCPAsZGIGjpK05BJPuv+0Vog1lfg4XpBMSZhXETYHgaMFDlc2YsRjmBA
I1oEA6NKJ37Hvnbv7Z7FKojtGLpkpg4ScxMZT8iMz7fOhSEOgQYLQy/afn5mDFwmvoxf8ta4w1wo
a2x6oMNcTnsFBnJ4c53EEZBopheuD+hQaoel3M2qA6nmKWy5KZgOifRhHI0M4qr3Pl4LuNee4Ohk
lwYHVBJm+sihxQCTx7GsyDbzP1A7ZKFF+AW3jiEwTf7y7SswvQd+FT3PEaqUOiN3ztcDvoiTq0Ud
AzX8BnniT+tYRNKuRc7e4g1qbNvSyFbJt9u2F45MoFFzyl1D0eAxgJbyKyiAPcXS7QEjGBHweFwn
GngCilKpOOizKRSDgrTWij3x0EhQCUYbUPBGw9lrhrLPO+C5U3rJv1oQtgmtYiQaMbDuxFQGqAui
ECOCERVrbit+vsZ40a9PEikZ4biodj6IiSMjALUCse6c/g+QTFLeg0CIfsGXVUqAe4OMCoOad+nC
/ATbNLniqtq+BweX9Hd4vMoHLMzeh85AwytjYcEOPRD1Mtyj4W83feAn8J8qzdtyqeasxsAq/XJm
OpGUGO6Kn2YcMHB8uChjxJA3ZSXJ5uKOMW0zA0ds/GF1XgabM0uVXdRhcHvIGwgwabpoiA/OWH2u
2EW2zzdvIllQ9oCvj3Ls7kWSTmgd4lDerp6FQq13LfiZIJBdOa0qph7NfrP+7n+sghDdQY536EgI
BqXlUROMO3XKd5e0GJW+ZAKh6Z+5xwJOLlQZr1/lootrj04kYlmQ4eO9KhXciATXC7xMtm8tiFco
vvboOkDfb3aA/mGAopAoZzNtduAtXwIpq0ZIaGy+cKVs3eSZ+yD8h+RPP4jlSNapCjedsoiC78ja
20vlv/AdZ7hgFqyVFZsJkyrgOWkuynU3IQmCoaRAUyka/m8FoxfrjOy6rio4Be/3OvThe3sgvIey
P38tT2aen4irvNWfMS+C9pgbax/F7TQUy8nBs8RlEUlRxKDEscWlkIbRrZlYj4oKzzo0KLM0GDfk
WPMi82Syfh2kb5r4GYobldM67jGVLdjgc1ZMkXRDmWKFDdXMVSYEFp5NYobZmQpv1EwoOCObg1gX
6DqoSN3f2OtQ6HN1sICE6CvMpJ+/axPefFcwV1zQB7K3l4W6yJlPIBrVPZXkPZFv7vZaorEteB6O
Gb2xHHC/OdN1G6Gg8naFksAl+d7RhbFk8TqUgbXK+V8gZOiHHfpZxVAzODFxjgxU1YLtEJKjTS4Q
sT8UFfKWCiMiQbokrEpHmzXw0nL5KBc7muZjxu+d/w8cwkTG1aheRnArLy7DH6nDMk3TCyRcT32S
i+tj6NpWCp5YLiKGGyTxr5T3yzZUTqhEDIBHy84aD9HJkFBuVz0TpU88sFfYY9yqybNIEHBE1jCu
GqPvv/qD9qFfwdObt1AlhyanRwkuMm+TDH0906/lQz6lvZ3MH9BERVb7+SfHLTB+5el6YKZWVjZO
ut5f8euUIV7g82xqc2XYwMUJZ7b+yj3m2lHPW6tMgulBVHUfnKxNkDo1FALdKA57B2VCqb5a5Wkr
ArMSjTTyLgzXnCTuO02426Cp9+eRelqiXF74fSH3Z/DFQlKlGWDWpo0xeE4O0gpL2pT+LSIw3SK7
93H8sj3Mc/wVJB45BMOzIPgVxJ41+l+AOgMbwyeKdWEQG+KaDrHBjchcmKh/jkuQui0qaL9UngrS
h1pELRa3I2iNucRC2FYSXxBl1Pv77+OXoQJ4rBTh+B62dQFAMiEd5Bc1GMo6DEc/laT97MoC+i2l
2Z8CBOibQmQ2bqX72K6vfAKFzabzGfk/VZWuFgpqoxnXm47DodNGo+bSjJZ4C1xZOinRHo22qbOx
wMVgt6NbJApRN3yIJEEAU74sW4Dvbo8gVMU1K0BNVNnuPu/toJDyk07c3Py0RiUihmO9xRVd4wXR
hNdrV+XTnzCwZrZ3dU8g7Cl8SLRWPy42ui3OuoRYkDPPTD2s2Y6pFG16zo0JdWd5dKno7E/eAd/q
ODyYuaC4L4mFCrjJNG4LUNeGa+CepmIVmWVLmnPLpIPFH7jL1Xiwov9thSnZoKtR98xb+jCqOISt
OIJKUQawXBsRoowe/Dxifgz73XTrrxenMj4EbvIPwHQ2D4bPGp4f4z4iaTzhObxmsP6/XZ7lWDiH
ArtoFijgcOEVfb0qweER/L4XZjL/0fDozHWL2qpO0BEiGl8cO3uhTSVe7acTgwXxCbw4DhgYQYOP
aVnqdnRsQ4venOpQp3XjpJAUQ4DuhylM0Yuu8lRsCYUfIEY7//KwfGIB9EbPooV1VOZh3wYrSJxv
23eQG8xCRZKIF+gS2g70YsyAwOd+/JNZSV5TJP/Nm43Qif4ZV3ZiM/Gzkekz7tRAi4jT7pu4Rp8k
bLBmXsgjPFDpjGkHIdctH6jceN702swJSq7a8N0pHPNTA2rw+k6DG+CAZyQnzzz6s5VagMp37A4w
qVgNwvBCR94KJBdnznshJNz7XFxRnj+fv3kq7vzbifEXtYMAdz7Vaej2lTIEmVd2Ccw6Wce80TDk
yfBrxi1SYclqbSFUbS2M+fS4JvTyR0tgp1chxCUFV/HP6IN77ODqazlC1Kcz9rpurKAUT1WdbrU7
/ZflnPYU1gzOeyoitqos4u4DQm+V1f6CnFOZ5RyYs33bpSOhsazuDRwtvuZAgrRFUDtiKQ/FBeKf
MRqkgPHrjLfp1FjaTWFvP0+AtSCxujQ1Qb+cl6bz+AXs1waouRd2P8eXUkChXasOmbejlqhQ3Jnq
XO+Abx54p84qXeUOR5IRzj/daYWhdQWzGw3XGRrmtX67oJfKmXjFWkGaRP95GkEYT3AkT5T+CEkM
2ZAcsZy1Ps4QrxEI45d5yz3pacfc2EYu0+MdBcfgi4UxJ0OTH9fXhSFo+Z+VD43LD6nIqyowTpSD
Jd6CBgG9v00uNmYtQ3f6q4nrjEDasYiIcJ+zKp3WiW7dCFmm3YtInMgzpuN/bp+2K8Vc+aourG8m
DhZAiRTYXOesBIaLZJpj5M6AOk4tNmMarG3gLVbHoaJA6MPMkkqL6z3/+6c3lJHbMWb6joDumjYi
FE5fvJbGMwmUcxjo6uNHpWi6ES4KM7Yk3o/y2yt9EeNFRMH1Ln5W42kBRC6XUtQl9z5HJYmRmyox
iVEJdkdBWIAWy6qKAf9UyOhBaN1aAaj+6gdLUP1TkgHUe9eoWNuxBk3bY7faxgyyDe+Gu2M7DgaC
GtUHMeQXMuHRH0HUr4JIAU5sAHB/Fy9/4PVSzq7I6si1NIsaleS9ZpQQ0PPvjXQxIqvLlJtgbTLp
qSaFUGVsc+mIHtcS+9Ah0B8t7/PX1EGUzeiIxCxGTxPTNrcbfX4Fu5FGNP+6pec18EKLKpGohrK2
TYGFm0WJGfgiUiajjY5dnnJtWmwMa/QGpg4OQlzmuD9JKahfdHzMi42vBplRWnU5DAWittU5wEX1
+FinJbol/oNY5Q15aDPVgHUrLrNNZVm9/nfSQjicwRurE/WmbQo7NAelYiJ8Iif1uiZeixxitLxV
axK0o1k9EJWc8pZa6tKoILCdXpfxVxeh2syevKd7v79Qt+S2hsJNQzMa4NctoQw+c6yjW/2VZmsl
nkkl1l4tmZloT1BRIv2idmrJQwRB3p/q3x+fSPTxkpkRlfxjQ8la3WAzxPul+7Dk6GKbi1cS1sJF
Azf865iB/ehpsrlIeLnwJREP0Q9DCO3iLwMJ3Ujgdt8KmWPgAHrGkj8YFU3Htw/S0tRobeHDPJlM
2rHpqE7RKaM6THu217733ZxbH/sxVrJhNcMJcgbf/XAfznFMwctK8pGmUwTNGQEocPwVKfLHne18
kL2ihT85vC2OEK/kDh20lJZzVQZIrStA3/O4rkk2IPnhp2k+e9L+lSnhdP833LX7btyIV5wTtIhK
yxxn51b87Not7kKSQwL81pmKsimFXowUl1K2Oo9QLUK0ZvW7irbHaXmAoa/b9kCjvoRIDcG24ZaA
/xeba2OVCXDkDyanwy1ERMkCdgmYxQaQa1uLRSEwWR+jT69RTIQ/HTvxnmFMnTER/0uduqacOqAG
bmTtT8Ua2eswhM9joSKCNGNKBHJL2fH1wXu8hEtdsHIch+XXhctKZsZqwK2chK8R1Tvd34tNwul1
ptHkYOWByhWtqZfzgDxiIONwmcwT3PctE5f/ZQeBYL1NyuhYh5TUo+qATCs7v0V5Vms1mnkLHSIb
Bu9zjUeCqy/jiSkdh0M1BSQCinN79xQXpWwjb4A+ed3jYnXu1QvQCwudIhbdR2s+DJZYJeP3kFnS
bUJm+25thlBsVaFxekteZrNfN4z1VGHfqUvM8azKBlPcHvEyTm5L7JVK+0C/U3BKcFQywwxyJwfS
TmLVE8tOLTZt2QRnuZnJLoK8klBTkBSsGQTAbQNt2wD8TIXZDCoeMDtsXtLCiWT5c5++RPd+HoO9
wF8zKWqwCHAFhWW5pILXPzYzkXFYE61WRYWJ/cz/s5u8LGvCPC/COaExfsDHH+AuWj90OXhJ3mNJ
pfJ0rFftT2lSrmadxCKePkMCGZ1nUJEQYv08dXXlmiJyDtWvvZEWGXE7ldWkfoK87hIHxqo8wKO0
FoOilLUGlwJmckqvjlkm6jbQZeF7sbsNda6C01HBekzCTUwHAFptr0uTpt/7Rv4uCDAsRxhZMVST
tLWTNJ+DDtj4BAZDdsmHAfWPl2sg8G3q7Uiwtt2o0JTKIcLg49qzfXU79Fc4aehL2pDwTF6UsYy/
42fU7sW8cfnelmMZ77YRBhhxIwbFqXYA7QOccPFwwz5hDPDKws6GT5AzhdqpM/TwGj818AGoClV+
UGNBQQMfnb5ft+Sj+OVRZ3cTU7R5bkuP0EoiSXh+88ec+phoWlL3x3qTIoyXDBT3xgg2V8OADB5y
/U+eaw5KoxA+5JX93swzDFouIu6MKLPPRDQv+bhemA1QPtNzs2Ez/mKaCoXsSd+NKb6B5WS9ib7+
De820Qk+/+amdetZHJp9fWjNdAIdrEHdxaAkzcVITP1C9S9XgXNNh6p9nqrJiQgk1TYoZJ+4Xbtq
027bcU8Sb7J0gZOroQJDdLH6ZqNjUZLEF326uImob3O/W+MidxZ2InlaMtD3/aIzFIJ4lYumtpkp
xq85lTQO234Rdv0ztApVivJ46C44+FVMsXgU3PDqptUsYvfzT0FiuQf2EqhgYplBxCDYUFM2wySM
kzaxwvyYNLFy9cPfj/9PaMJ1waJ1JicOnBrYWZSXQr/6f/5Bn24dUuQF//UOylwfPZO69tuGVKOT
ZGdkE852kHp8pR+XFT6jRZXAuVd17BFsPNpmE+MhbQaImiRNMf0Bcw/ARKT7wt+qGXaQsRp4CiwD
6IHkiEsM1tP5enVgw4JEt74mJp6zSo+JRHzmLNYXVIWZckOzwhWMbnQhNuCaRUv8zw5vOGidnjQM
VBS9U2kiwdsKjhX+w9iwEUkYHhxcCQOlgXIj6BT8hxaqNZjN2R4hnRUbLpgUFByroFtzcMKskMXy
surfXZYfeo5n/GvZzDO8MY1eow8KSmKG2rZ0uRQJiuXEHa74f9cKbwMzpeC42pzNZhX1j1l1zpIP
8Kv8ezB97Q86bGy4J1681dpms/2XtAHNNvpi57eonw9rChDcteBYViPCT6u2JDyJaVfE+H4T+BAy
4+jWYETaSiz8vXmFUaEp/mfubIpJ0v+sS/UT5ejs5WBvfmMzveOJCA7xN5wY3qaTMtOv2Ubi4K8T
xupAubefnyAoALtfqnLv6bstLEggRQn28xFm0ZM/SFxK2efjLB0nB/kDb00rkTYDZRsgpYREqy6D
X6XwZ5rTayU41S5Q3TbdyGv84/TpQJ38eaQTDc381aljLK8O4LZ7GeWnGDbexoGMtEUD+ohb2SjC
0SZaOvXfyj9pmiUfmZ4tbWUfaayf5mGJPleg1SO3/66EtpEJYZq/51B06hOGJweI9lPuLtD/6ZbO
8iOV3SLYToLYvgX2tB0F7MbCc4BwgZz+J2pkzJMyBUgFgHJAPtCIk5K4sQe8mk+dgBThiPZEdV0h
Jd6rk0JUNNSd5ZxGACfE3C055/Atz2KFuMH1QW2SsnT9nYwvlABBvX31lrA777J5eZVQVhc1QJmr
+BgFcPzmpFRvK0F1ilc7AZohKk2GdeulKmYhofJe+tudwvpRMuXQ3wht5tNByDRerktfN+v6OP88
MsWZk3arngU2OIJS7LpjEER+rv9lyBdaNecv+M+PoKo91vk/qc1kP3pz33G2o1SY+md501wlMW3P
Uz3We+Ka1cWYOnIVgEH5tXAn1nuXSeM4veaunhBX5+kOTp578+zMh9wKFkxEAdCMgxPRfwhvvroU
blOXfLbfaddENhGx/qPa7kJ2dIx/H5+h7oqelWFYQdLmR+r0KR2w4oFb/N3dfSyrwe9P7H6k7Cle
r3IEhgcVycZil1Qv82dQ4CdUh9iuDuBsS1eRP5rbERsXA11lufGK+h0ny19iJtknz2aJ2iDz6cDu
dlbEIJoJLojG7mrcIAuHGUwvswuK6P+fR1FS+orvWW8YAOS1ri0RLVezTSIAZ6FHC+WG6SgLkjc/
kfLpnEp7Kl+QUHxpmJRbFNzDd+AMYIX9976AU2qpmIU/IpeXe9L9eh+REQhh4oV8UNgUIa+/CetG
UiLLvj3J/lAhh0T6+iyhhxXB5AzYksLKuY0/RrLlUzTHDBX1ejQ4qJoynvgoZp0ZBo/FBCMbWg5V
oztrPPH25Ue460lPQ8h3Lg8peV7MJ2r89tO2i2RsepsXLxYyWc1y8YlQPGhxm4hk+n9R9KlCLCBB
jLTd3zKVmZDqbywnKDhUnhtOHQIBBamS6Obhs3Nv+OFTaxo1oZq5+Jb624Vn3v8xaGCg+wduXUTk
OAkIVn8olLIDZNk+Mm5h35ZAse/MciA1X9OGwqfGafKE1UrrMb/LivWKPNk+M0byYbC117vmqYsF
14xu8vF94sdSFeieVaq+ulwkXNGN9htpnTh00Lg7is54M6onv3q7lIy05vgnyTCDZ+RK5WUR83sK
fpMIs+1cnCwvSTibzrW6NycrlKy+xZfU2RJdTDi6nkEO6T1qc7ItDu+3+5xDqhfJ9s1rQfh+v4Gj
i/Q3lXS+ABuUWtbLUDcf8n874Mw0aqzYsCnLV3G9z9wT3Fwl82uxbHKwISd8CAmnOmm6JF4lgKP+
q3NUXQFMvoSNhqejrIGAVkAtL+Qp5LnW6h4i2GHeNXBFY0iYfHZHsPUzEFOcwFjM+LgBkOx4LmJ3
XB9UX2jNNPy5WbRbuXWsIH8lEuyA+39XHLzp5nw7bLPN6bgO5mBmYZ1Jyb7XHRQg+KR68pP8eHMe
olXcFGC77jeJOzx8yImJZdBrYyNtmcyeDYZrwoxqp+fXHc/zyT2vG9lmmvoaPImTKgXHFCg/Ew3u
CV+DdlF7Eu+HgNxdPhti0Nnd81inh5NkjtJyy5Q6Yh2qLK8aBjn9HGUx0x35dKyr08HXJDXX9pBE
weBErWHCVazpST3oVOS2g8qjboG/LTo2Sws9q6vqYSPP93+fDM7t5JzzcPwLdok+GVg50a+0+lNS
cDpAA+Qp4Pqn/WBIqqB9rOujBq6PSRfCBAkICbzG/q5oc76eFf5iL9XRgWjYSOlLOQ5uTBeJPB6v
Na02fRniQ+IY1veiokf+BrbTjtBrHJhxny2ShHD8iTPtnujB4NPQodROtwu8/LhUwQv51+fsolt1
hWqHrOeTmSn5efp7Ku+ONUkRns/BgWlF+ZoDK2F9LaXBpJ6HGW+PaLikiNfO+su8deUd4+Q0wFlY
TwDQXFr8Y1UXIX1xKH/81nqijQVugYv0a9H/t6S9ieZBzImj72ljHrN0Rm40HrZY6IR3WNO3puop
RfKfEFjDLiebr9YfdYsk16x40judX7x9UKU9GQuXU1X+35u4lhQWLJHrTdIBWbWY2ciugORh8lg0
2To+tv7+HmzbL2tZ8vi1fHfqOUlKbqHe5Z92IaId2l5klbgRgA8VLp/YN7s3YUBiroPpQ+ifcUjS
1zThKfKf74ENCco2lyU60zx7FHImzAfSCjrFM82mmhtlojZ3Fn2CR2HhvHQcEWy9Z1Q0H8OIgFRx
czYQ/wtjR283RCTQGecHUuYfXnlY8BwVc0qI9JUtJxBYjnPzaoEZP4mLUE4DjAzYn+3C6a6xaszV
jsqWKfMU7Pd9BR9OAu55ammlAyej9a6S6rNG9WDCekSqeH1VEJ91mSRRwkUwsl5C6GetMd47yy3Y
RYH0lWzNZbRYRhRWjRDg2/jsSOv/l/081D/Fn/yiPMFDT/TFG+XoDAJU4uqW4sngeIG8ozuaCfkQ
X3w1OuNhWngLBawPNA1QuLMiqQ32Nw1ytJwVTQs0TMeo/ONaUOjIHJz4pv8w30JCFBu3qwvnLItK
XAtujqLlo1S2x6YYMXI8nY+MF4tBUD3T7S8F8lTy9Pi3MTEas3xEaYJd5VlKW7sv6Y5fRqHTV8vt
QqolMgiHa3Y07ozc4jmYMdbH62Ll+DBnlmfrBfw2JAlZYXNq0dsm7Ft9H2otlO+FVSG8gKsu9Dfe
T0ZdiMnvkSDePFvydK9AyjyN33CwBaVkfCpvSfHGUGdFkmdM5XUuIy0zxu7tz7wOR2vECHPgNQus
cjG1LT3SfJmDkg+JIvmQGcJhjpHvbBAfr773kLYE9cHyjNUrfahg2GOXneXy9Faf8oegmEwhz0Ct
yx6OhKSkAgACXOw1DK59AxNgXXvt9k+h5k+vmDXbGHbGJN4e2TTHoA+p7UZ+gTY2pnPylytzez6O
JG5soUDG3EXbsMq3ixn/BOeRZot1stNefFBE4F51xuY3kyMi6GTKTR7CWpF72BHdzI0f2TIjT0lA
tfX83Nf7LwzHULx/vgbVFEYzv1GBBgrA20R6p/JuYtzhC5wp+1vJuTdauBN74CkEWKvCsU6DlDb9
Pygo8b4R1Ny7IRrq9B7UrWAZ0MHppa8WZ/TVUOJoQ4Z87YK6ziTzBIGea7+zCdhuch/B2qcyqnCu
fsJDY5ium5poBamwJXEP2w1pKi9bbnuUpvTV2KfCYVqGA6fa4CwvcA/O4x7i52L1CZfd/Q1wPzeH
0MO2BpiGwH/jPgAuehCNmL4tBsVSLSlCcBsxOPwF9qegcba+Mn7+6CB3B2vKXAB2C3hXO64+RO79
XV37/qbNIl3FSlYbrKGX3GRR1YLIGYpPo3lkTCBp06vCwtD4rKVPjk9/vdh3c0gFzBd7YNRho6CC
dNqU91vL+AEji6DXmyQoSYnUbIt/Y/g5BQ3s3s2qwn7URCouCS6olxmQC0GuRQgZYXxV+QgTvysb
az/HKb2uc/5MDQTvv/2LjYmGjddTOf9BZDGqzQ+xvVq8TLO8tPusLASABSVWff08vesfSn1s2NR8
b/XuNcTw6mbRINHLF5mLyDsy4dI1OmhNxWobfxeR8upFvedmVbZdCpa+wqU1JCVw51DFPV2nhsEg
UlDG2Xr7YpGH
`protect end_protected
